../../src/verilog/alu.sv