../../src/verilog/multiplier.sv