../../src/verilog/mux8x1.sv