library verilog;
use verilog.vl_types.all;
entity mux32x1_testbench is
end mux32x1_testbench;
