../../src/verilog/mux4x1.sv