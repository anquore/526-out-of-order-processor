library verilog;
use verilog.vl_types.all;
entity decoder2x4_testbench is
end decoder2x4_testbench;
