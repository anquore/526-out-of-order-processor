../../src/verilog/mux2x64.sv