module multiplier(out, valid_out, A, B, valid_in, reset, clk);
	output [63:0] out;
	output valid_out;
	input [63:0] A, B;
	input valid_in, clk, reset;
	
	//timing module and register, 4 cycle process
	wire [63:0] Ar, Br;
	wire v1, v2, v3, v4;
	registerX64 regA(.out(Ar[63:0]), .in(A[63:0]), .rst(reset), .clk(v1));
	registerX64 regB(.out(Br[63:0]), .in(B[63:0]), .rst(reset), .clk(v1));
	D_FF valid0(.q(v1), .d(valid_in), .reset(reset), .clk);
	D_FF valid1(.q(v2), .d(v1), .reset(reset), .clk);
	D_FF valid2(.q(v3), .d(v2), .reset(reset), .clk);
	D_FF valid3(.q(v4), .d(v3), .reset(reset), .clk(clk&(v3|v2|v1)));
	assign valid_out = v4&(~((v2&~v3)|(v1&~v2)));
	
	wire [63:0][63:0] ands;
	wire [62:0][62:0] addeds;
	wire [62:0][62:0] carries;
	
		andifier a7(.outs(ands[7][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[7]}}));
	andifier a6(.outs(ands[6][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[6]}}));
	andifier a5(.outs(ands[5][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[5]}}));
	andifier a4(.outs(ands[4][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[4]}}));
	andifier a3(.outs(ands[3][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[3]}}));
	andifier a2(.outs(ands[2][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[2]}}));
	andifier a1(.outs(ands[1][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[1]}}));
	andifier a0(.outs(ands[0][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[0]}}));
		andifier a15(.outs(ands[15][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[15]}}));
	andifier a14(.outs(ands[14][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[14]}}));
	andifier a13(.outs(ands[13][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[13]}}));
	andifier a12(.outs(ands[12][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[12]}}));
	andifier a11(.outs(ands[11][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[11]}}));
	andifier a10(.outs(ands[10][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[10]}}));
	andifier a9(.outs(ands[9][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[9]}}));
	andifier a8(.outs(ands[8][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[8]}}));
		andifier a23(.outs(ands[23][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[23]}}));
	andifier a22(.outs(ands[22][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[22]}}));
	andifier a21(.outs(ands[21][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[21]}}));
	andifier a20(.outs(ands[20][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[20]}}));
	andifier a19(.outs(ands[19][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[19]}}));
	andifier a18(.outs(ands[18][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[18]}}));
	andifier a17(.outs(ands[17][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[17]}}));
	andifier a16(.outs(ands[16][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[16]}}));
		andifier a31(.outs(ands[31][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[31]}}));
	andifier a30(.outs(ands[30][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[30]}}));
	andifier a29(.outs(ands[29][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[29]}}));
	andifier a28(.outs(ands[28][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[28]}}));
	andifier a27(.outs(ands[27][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[27]}}));
	andifier a26(.outs(ands[26][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[26]}}));
	andifier a25(.outs(ands[25][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[25]}}));
	andifier a24(.outs(ands[24][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[24]}}));
		andifier a39(.outs(ands[39][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[39]}}));
	andifier a38(.outs(ands[38][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[38]}}));
	andifier a37(.outs(ands[37][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[37]}}));
	andifier a36(.outs(ands[36][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[36]}}));
	andifier a35(.outs(ands[35][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[35]}}));
	andifier a34(.outs(ands[34][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[34]}}));
	andifier a33(.outs(ands[33][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[33]}}));
	andifier a32(.outs(ands[32][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[32]}}));
		andifier a47(.outs(ands[47][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[47]}}));
	andifier a46(.outs(ands[46][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[46]}}));
	andifier a45(.outs(ands[45][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[45]}}));
	andifier a44(.outs(ands[44][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[44]}}));
	andifier a43(.outs(ands[43][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[43]}}));
	andifier a42(.outs(ands[42][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[42]}}));
	andifier a41(.outs(ands[41][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[41]}}));
	andifier a40(.outs(ands[40][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[40]}}));
		andifier a55(.outs(ands[55][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[55]}}));
	andifier a54(.outs(ands[54][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[54]}}));
	andifier a53(.outs(ands[53][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[53]}}));
	andifier a52(.outs(ands[52][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[52]}}));
	andifier a51(.outs(ands[51][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[51]}}));
	andifier a50(.outs(ands[50][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[50]}}));
	andifier a49(.outs(ands[49][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[49]}}));
	andifier a48(.outs(ands[48][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[48]}}));
		andifier a63(.outs(ands[63][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[63]}}));
	andifier a62(.outs(ands[62][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[62]}}));
	andifier a61(.outs(ands[61][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[61]}}));
	andifier a60(.outs(ands[60][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[60]}}));
	andifier a59(.outs(ands[59][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[59]}}));
	andifier a58(.outs(ands[58][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[58]}}));
	andifier a57(.outs(ands[57][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[57]}}));
	andifier a56(.outs(ands[56][63:0]), .ins1(Ar[63:0]), .ins0({64{Br[56]}}));
	
	//full adders
		assign out[0]=ands[0][0];
	fullAdderArray63 line0(.S(addeds[0][62:0]), .Cout(carries[0][62:0]), .A(ands[1][62:0]), .B({~ands[0][63], ands[0][62:1]}), .Cin({63{1'b0}}));
	assign out[1]=addeds[0][0];
	fullAdderArray63 line1(.S(addeds[1][62:0]), .Cout(carries[1][62:0]), .A({~ands[1][63], addeds[0][62:1]}), .B(ands[2][62:0]), .Cin(carries[0][62:0]));
	assign out[2]=addeds[1][0];
	fullAdderArray63 line2(.S(addeds[2][62:0]), .Cout(carries[2][62:0]), .A({~ands[2][63], addeds[1][62:1]}), .B(ands[3][62:0]), .Cin(carries[1][62:0]));
	assign out[3]=addeds[2][0];
	fullAdderArray63 line3(.S(addeds[3][62:0]), .Cout(carries[3][62:0]), .A({~ands[3][63], addeds[2][62:1]}), .B(ands[4][62:0]), .Cin(carries[2][62:0]));
	assign out[4]=addeds[3][0];
	fullAdderArray63 line4(.S(addeds[4][62:0]), .Cout(carries[4][62:0]), .A({~ands[4][63], addeds[3][62:1]}), .B(ands[5][62:0]), .Cin(carries[3][62:0]));
	assign out[5]=addeds[4][0];
	fullAdderArray63 line5(.S(addeds[5][62:0]), .Cout(carries[5][62:0]), .A({~ands[5][63], addeds[4][62:1]}), .B(ands[6][62:0]), .Cin(carries[4][62:0]));
	assign out[6]=addeds[5][0];
	fullAdderArray63 line6(.S(addeds[6][62:0]), .Cout(carries[6][62:0]), .A({~ands[6][63], addeds[5][62:1]}), .B(ands[7][62:0]), .Cin(carries[5][62:0]));
	assign out[7]=addeds[6][0];
		fullAdderArray63 line7(.S(addeds[7][62:0]), .Cout(carries[7][62:0]), .A({~ands[7][63], addeds[6][62:1]}), .B(ands[8][62:0]), .Cin(carries[6][62:0]));
		assign out[8]=addeds[7][0];
	fullAdderArray63 line8(.S(addeds[8][62:0]), .Cout(carries[8][62:0]), .A({~ands[8][63], addeds[7][62:1]}), .B(ands[9][62:0]), .Cin(carries[7][62:0]));
	assign out[9]=addeds[8][0];
	fullAdderArray63 line9(.S(addeds[9][62:0]), .Cout(carries[9][62:0]), .A({~ands[9][63], addeds[8][62:1]}), .B(ands[10][62:0]), .Cin(carries[8][62:0]));
	assign out[10]=addeds[9][0];
	fullAdderArray63 line10(.S(addeds[10][62:0]), .Cout(carries[10][62:0]), .A({~ands[10][63], addeds[9][62:1]}), .B(ands[11][62:0]), .Cin(carries[9][62:0]));
	assign out[11]=addeds[10][0];
	fullAdderArray63 line11(.S(addeds[11][62:0]), .Cout(carries[11][62:0]), .A({~ands[11][63], addeds[10][62:1]}), .B(ands[12][62:0]), .Cin(carries[10][62:0]));
	assign out[12]=addeds[11][0];
	fullAdderArray63 line12(.S(addeds[12][62:0]), .Cout(carries[12][62:0]), .A({~ands[12][63], addeds[11][62:1]}), .B(ands[13][62:0]), .Cin(carries[11][62:0]));
	assign out[13]=addeds[12][0];
	fullAdderArray63 line13(.S(addeds[13][62:0]), .Cout(carries[13][62:0]), .A({~ands[13][63], addeds[12][62:1]}), .B(ands[14][62:0]), .Cin(carries[12][62:0]));
	assign out[14]=addeds[13][0];
	fullAdderArray63 line14(.S(addeds[14][62:0]), .Cout(carries[14][62:0]), .A({~ands[14][63], addeds[13][62:1]}), .B(ands[15][62:0]), .Cin(carries[13][62:0]));
	assign out[15]=addeds[14][0];
	fullAdderArray63 line15(.S(addeds[15][62:0]), .Cout(carries[15][62:0]), .A({~ands[15][63], addeds[14][62:1]}), .B(ands[16][62:0]), .Cin(carries[14][62:0]));
	assign out[16]=addeds[15][0];
	fullAdderArray63 line16(.S(addeds[16][62:0]), .Cout(carries[16][62:0]), .A({~ands[16][63], addeds[15][62:1]}), .B(ands[17][62:0]), .Cin(carries[15][62:0]));
	assign out[17]=addeds[16][0];
	fullAdderArray63 line17(.S(addeds[17][62:0]), .Cout(carries[17][62:0]), .A({~ands[17][63], addeds[16][62:1]}), .B(ands[18][62:0]), .Cin(carries[16][62:0]));
	assign out[18]=addeds[17][0];
	fullAdderArray63 line18(.S(addeds[18][62:0]), .Cout(carries[18][62:0]), .A({~ands[18][63], addeds[17][62:1]}), .B(ands[19][62:0]), .Cin(carries[17][62:0]));
	assign out[19]=addeds[18][0];
	fullAdderArray63 line19(.S(addeds[19][62:0]), .Cout(carries[19][62:0]), .A({~ands[19][63], addeds[18][62:1]}), .B(ands[20][62:0]), .Cin(carries[18][62:0]));
	assign out[20]=addeds[19][0];
	fullAdderArray63 line20(.S(addeds[20][62:0]), .Cout(carries[20][62:0]), .A({~ands[20][63], addeds[19][62:1]}), .B(ands[21][62:0]), .Cin(carries[19][62:0]));
	assign out[21]=addeds[20][0];
	fullAdderArray63 line21(.S(addeds[21][62:0]), .Cout(carries[21][62:0]), .A({~ands[21][63], addeds[20][62:1]}), .B(ands[22][62:0]), .Cin(carries[20][62:0]));
	assign out[22]=addeds[21][0];
	fullAdderArray63 line22(.S(addeds[22][62:0]), .Cout(carries[22][62:0]), .A({~ands[22][63], addeds[21][62:1]}), .B(ands[23][62:0]), .Cin(carries[21][62:0]));
	assign out[23]=addeds[22][0];
	fullAdderArray63 line23(.S(addeds[23][62:0]), .Cout(carries[23][62:0]), .A({~ands[23][63], addeds[22][62:1]}), .B(ands[24][62:0]), .Cin(carries[22][62:0]));
	assign out[24]=addeds[23][0];
	fullAdderArray63 line24(.S(addeds[24][62:0]), .Cout(carries[24][62:0]), .A({~ands[24][63], addeds[23][62:1]}), .B(ands[25][62:0]), .Cin(carries[23][62:0]));
	assign out[25]=addeds[24][0];
	fullAdderArray63 line25(.S(addeds[25][62:0]), .Cout(carries[25][62:0]), .A({~ands[25][63], addeds[24][62:1]}), .B(ands[26][62:0]), .Cin(carries[24][62:0]));
	assign out[26]=addeds[25][0];
	fullAdderArray63 line26(.S(addeds[26][62:0]), .Cout(carries[26][62:0]), .A({~ands[26][63], addeds[25][62:1]}), .B(ands[27][62:0]), .Cin(carries[25][62:0]));
	assign out[27]=addeds[26][0];
	fullAdderArray63 line27(.S(addeds[27][62:0]), .Cout(carries[27][62:0]), .A({~ands[27][63], addeds[26][62:1]}), .B(ands[28][62:0]), .Cin(carries[26][62:0]));
	assign out[28]=addeds[27][0];
	fullAdderArray63 line28(.S(addeds[28][62:0]), .Cout(carries[28][62:0]), .A({~ands[28][63], addeds[27][62:1]}), .B(ands[29][62:0]), .Cin(carries[27][62:0]));
	assign out[29]=addeds[28][0];
	fullAdderArray63 line29(.S(addeds[29][62:0]), .Cout(carries[29][62:0]), .A({~ands[29][63], addeds[28][62:1]}), .B(ands[30][62:0]), .Cin(carries[28][62:0]));
	assign out[30]=addeds[29][0];
	fullAdderArray63 line30(.S(addeds[30][62:0]), .Cout(carries[30][62:0]), .A({~ands[30][63], addeds[29][62:1]}), .B(ands[31][62:0]), .Cin(carries[29][62:0]));
	assign out[31]=addeds[30][0];
	fullAdderArray63 line31(.S(addeds[31][62:0]), .Cout(carries[31][62:0]), .A({~ands[31][63], addeds[30][62:1]}), .B(ands[32][62:0]), .Cin(carries[30][62:0]));
	assign out[32]=addeds[31][0];
	fullAdderArray63 line32(.S(addeds[32][62:0]), .Cout(carries[32][62:0]), .A({~ands[32][63], addeds[31][62:1]}), .B(ands[33][62:0]), .Cin(carries[31][62:0]));
	assign out[33]=addeds[32][0];
	fullAdderArray63 line33(.S(addeds[33][62:0]), .Cout(carries[33][62:0]), .A({~ands[33][63], addeds[32][62:1]}), .B(ands[34][62:0]), .Cin(carries[32][62:0]));
	assign out[34]=addeds[33][0];
	fullAdderArray63 line34(.S(addeds[34][62:0]), .Cout(carries[34][62:0]), .A({~ands[34][63], addeds[33][62:1]}), .B(ands[35][62:0]), .Cin(carries[33][62:0]));
	assign out[35]=addeds[34][0];
	fullAdderArray63 line35(.S(addeds[35][62:0]), .Cout(carries[35][62:0]), .A({~ands[35][63], addeds[34][62:1]}), .B(ands[36][62:0]), .Cin(carries[34][62:0]));
	assign out[36]=addeds[35][0];
	fullAdderArray63 line36(.S(addeds[36][62:0]), .Cout(carries[36][62:0]), .A({~ands[36][63], addeds[35][62:1]}), .B(ands[37][62:0]), .Cin(carries[35][62:0]));
	assign out[37]=addeds[36][0];
	fullAdderArray63 line37(.S(addeds[37][62:0]), .Cout(carries[37][62:0]), .A({~ands[37][63], addeds[36][62:1]}), .B(ands[38][62:0]), .Cin(carries[36][62:0]));
	assign out[38]=addeds[37][0];
	fullAdderArray63 line38(.S(addeds[38][62:0]), .Cout(carries[38][62:0]), .A({~ands[38][63], addeds[37][62:1]}), .B(ands[39][62:0]), .Cin(carries[37][62:0]));
	assign out[39]=addeds[38][0];
	fullAdderArray63 line39(.S(addeds[39][62:0]), .Cout(carries[39][62:0]), .A({~ands[39][63], addeds[38][62:1]}), .B(ands[40][62:0]), .Cin(carries[38][62:0]));
	assign out[40]=addeds[39][0];
	fullAdderArray63 line40(.S(addeds[40][62:0]), .Cout(carries[40][62:0]), .A({~ands[40][63], addeds[39][62:1]}), .B(ands[41][62:0]), .Cin(carries[39][62:0]));
	assign out[41]=addeds[40][0];
	fullAdderArray63 line41(.S(addeds[41][62:0]), .Cout(carries[41][62:0]), .A({~ands[41][63], addeds[40][62:1]}), .B(ands[42][62:0]), .Cin(carries[40][62:0]));
	assign out[42]=addeds[41][0];
	fullAdderArray63 line42(.S(addeds[42][62:0]), .Cout(carries[42][62:0]), .A({~ands[42][63], addeds[41][62:1]}), .B(ands[43][62:0]), .Cin(carries[41][62:0]));
	assign out[43]=addeds[42][0];
	fullAdderArray63 line43(.S(addeds[43][62:0]), .Cout(carries[43][62:0]), .A({~ands[43][63], addeds[42][62:1]}), .B(ands[44][62:0]), .Cin(carries[42][62:0]));
	assign out[44]=addeds[43][0];
	fullAdderArray63 line44(.S(addeds[44][62:0]), .Cout(carries[44][62:0]), .A({~ands[44][63], addeds[43][62:1]}), .B(ands[45][62:0]), .Cin(carries[43][62:0]));
	assign out[45]=addeds[44][0];
	fullAdderArray63 line45(.S(addeds[45][62:0]), .Cout(carries[45][62:0]), .A({~ands[45][63], addeds[44][62:1]}), .B(ands[46][62:0]), .Cin(carries[44][62:0]));
	assign out[46]=addeds[45][0];
	fullAdderArray63 line46(.S(addeds[46][62:0]), .Cout(carries[46][62:0]), .A({~ands[46][63], addeds[45][62:1]}), .B(ands[47][62:0]), .Cin(carries[45][62:0]));
	assign out[47]=addeds[46][0];
	fullAdderArray63 line47(.S(addeds[47][62:0]), .Cout(carries[47][62:0]), .A({~ands[47][63], addeds[46][62:1]}), .B(ands[48][62:0]), .Cin(carries[46][62:0]));
	assign out[48]=addeds[47][0];
	fullAdderArray63 line48(.S(addeds[48][62:0]), .Cout(carries[48][62:0]), .A({~ands[48][63], addeds[47][62:1]}), .B(ands[49][62:0]), .Cin(carries[47][62:0]));
	assign out[49]=addeds[48][0];
	fullAdderArray63 line49(.S(addeds[49][62:0]), .Cout(carries[49][62:0]), .A({~ands[49][63], addeds[48][62:1]}), .B(ands[50][62:0]), .Cin(carries[48][62:0]));
	assign out[50]=addeds[49][0];
	fullAdderArray63 line50(.S(addeds[50][62:0]), .Cout(carries[50][62:0]), .A({~ands[50][63], addeds[49][62:1]}), .B(ands[51][62:0]), .Cin(carries[49][62:0]));
	assign out[51]=addeds[50][0];
	fullAdderArray63 line51(.S(addeds[51][62:0]), .Cout(carries[51][62:0]), .A({~ands[51][63], addeds[50][62:1]}), .B(ands[52][62:0]), .Cin(carries[50][62:0]));
	assign out[52]=addeds[51][0];
	fullAdderArray63 line52(.S(addeds[52][62:0]), .Cout(carries[52][62:0]), .A({~ands[52][63], addeds[51][62:1]}), .B(ands[53][62:0]), .Cin(carries[51][62:0]));
	assign out[53]=addeds[52][0];
	fullAdderArray63 line53(.S(addeds[53][62:0]), .Cout(carries[53][62:0]), .A({~ands[53][63], addeds[52][62:1]}), .B(ands[54][62:0]), .Cin(carries[52][62:0]));
	assign out[54]=addeds[53][0];
	fullAdderArray63 line54(.S(addeds[54][62:0]), .Cout(carries[54][62:0]), .A({~ands[54][63], addeds[53][62:1]}), .B(ands[55][62:0]), .Cin(carries[53][62:0]));
	assign out[55]=addeds[54][0];
	fullAdderArray63 line55(.S(addeds[55][62:0]), .Cout(carries[55][62:0]), .A({~ands[55][63], addeds[54][62:1]}), .B(ands[56][62:0]), .Cin(carries[54][62:0]));
	assign out[56]=addeds[55][0];
	fullAdderArray63 line56(.S(addeds[56][62:0]), .Cout(carries[56][62:0]), .A({~ands[56][63], addeds[55][62:1]}), .B(ands[57][62:0]), .Cin(carries[55][62:0]));
	assign out[57]=addeds[56][0];
	fullAdderArray63 line57(.S(addeds[57][62:0]), .Cout(carries[57][62:0]), .A({~ands[57][63], addeds[56][62:1]}), .B(ands[58][62:0]), .Cin(carries[56][62:0]));
	assign out[58]=addeds[57][0];
	fullAdderArray63 line58(.S(addeds[58][62:0]), .Cout(carries[58][62:0]), .A({~ands[58][63], addeds[57][62:1]}), .B(ands[59][62:0]), .Cin(carries[57][62:0]));
	assign out[59]=addeds[58][0];
	fullAdderArray63 line59(.S(addeds[59][62:0]), .Cout(carries[59][62:0]), .A({~ands[59][63], addeds[58][62:1]}), .B(ands[60][62:0]), .Cin(carries[58][62:0]));
	assign out[60]=addeds[59][0];
	fullAdderArray63 line60(.S(addeds[60][62:0]), .Cout(carries[60][62:0]), .A({~ands[60][63], addeds[59][62:1]}), .B(ands[61][62:0]), .Cin(carries[59][62:0]));
	assign out[61]=addeds[60][0];
	fullAdderArray63 line61(.S(addeds[61][62:0]), .Cout(carries[61][62:0]), .A({~ands[61][63], addeds[60][62:1]}), .B(ands[62][62:0]), .Cin(carries[60][62:0]));
	assign out[62]=addeds[61][0];
	fullAdderArray63 line62(.S(addeds[62][62:0]), .Cout(carries[62][62:0]), .A({~ands[62][63], addeds[61][62:1]}), .B(~ands[63][62:0]), .Cin(carries[61][62:0]));
	assign out[63]=addeds[62][0];
endmodule

module multiplier_testbench;
	wire [63:0] out;
	wire valid_out;
	reg [63:0] A, B;
	reg valid_in, clk;
	multiplier DUT(.out, .valid_out, .A, .B, .valid_in, .clk);
	
	initial begin
	valid_in=0; //purely combinational test, ignoring valid_out cycle counter and clock
	clk=0;
	A = 64'h0000_0000_0000_0000;
	B = 64'h0000_0000_0000_0000;
	valid_in=1;	#5;	clk=1;	#5;	clk=0;	valid_in=0;	#5;	clk=1;	#5;	clk=0;	#5;
	A = 64'h0000_0000_00A0_FFFF;
	B = 64'h0000_0000_0000_0000;
	valid_in=1;	#5;	clk=1;	#5;	clk=0;	valid_in=0;	#5;	clk=1;	#5;	clk=0;	#5;
	A = 64'h0000_0000_0000_0001;
	B = 64'h0000_0000_0000_0001;
	valid_in=1;	#5;	clk=1;	#5;	clk=0;	valid_in=0;	#5;	clk=1;	#5;	clk=0;	#5;
	A = 64'h0000_0000_0000_0002;
	B = 64'h0000_0000_0000_0001;
	valid_in=1;	#5;	clk=1;	#5;	clk=0;	valid_in=0;	#5;	clk=1;	#5;	clk=0;	#5;
	A = 64'h0000_0000_0000_0001;
	B = 64'h0000_0000_0000_0002;
	valid_in=1;	#5;	clk=1;	#5;	clk=0;	valid_in=0;	#5;	clk=1;	#5;	clk=0;	#5;
	A = 64'h0000_0000_0000_0010;
	B = 64'h0000_0000_0000_0010;
	valid_in=1;	#5;	clk=1;	#5;	clk=0;	valid_in=0;	#5;	clk=1;	#5;	clk=0;	#5;
	A = 64'h0F02_0400_0654_1323;
	B = 64'h0000_0000_0000_0002;
	valid_in=1;	#5;	clk=1;	#5;	clk=0;	valid_in=0;	#5;	clk=1;	#5;	clk=0;	#5;
	A = 64'h0F02_0400_1454_1323;
	B = 64'h0000_0000_0000_0003;
	valid_in=1;	#5;	clk=1;	#5;	clk=0;	valid_in=0;	#5;	clk=1;	#5;	clk=0;	#5;
	A = 64'h0000_0000_5F72_AA7D;
	B = 64'h0000_0000_F29B_CF54;
	valid_in=1;	#5;	clk=1;	#5;	clk=0;	valid_in=0;	#5;	clk=1;	#5;	clk=0;	#5;
	A = 64'hFFFF_FFFF_FFFF_FFFF;
	B = 64'hFFFF_FFFF_FFFF_FFFF;
	valid_in=1;	#5;	clk=1;	#5;	clk=0;	valid_in=0;	#5;	clk=1;	#5;	clk=0;	#5;
	A = 64'h0000_0000_0000_0001;
	B = 64'hFFFF_FFFF_FFFF_FFFF;
	valid_in=1;	#5;	clk=1;	#5;	clk=0;	valid_in=0;	#5;	clk=1;	#5;	clk=0;	#5;
	A = 64'hFFFF_FFFF_FFFF_FFFF;
	B = 64'h0000_0000_0000_0001;
	valid_in=1;	#5;	clk=1;	#5;	clk=0;	valid_in=0;	#5;	clk=1;	#5;	clk=0;	#5;
	A = 64'h529A_8CE2_59F5_3AB9;
	B = 64'hFFFF_FFFF_FFFF_FFFF;
	#5;	valid_in=1;	#5;	clk=1;	#5;	clk=0; //testing valid_out (using the clock)
	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	valid_in=0;	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	valid_in=1;	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	valid_in=0;
	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	valid_in=1;
	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	#5;	clk=1;	#5;	clk=0;
	end
endmodule
