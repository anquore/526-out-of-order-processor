../../src/verilog/regReadAndWriteStage.sv