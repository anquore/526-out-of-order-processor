library verilog;
use verilog.vl_types.all;
entity mux16x1_testbench is
end mux16x1_testbench;
