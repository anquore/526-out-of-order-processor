../../src/verilog/mux32x1.sv