library verilog;
use verilog.vl_types.all;
entity signExtend26_testbench is
end signExtend26_testbench;
