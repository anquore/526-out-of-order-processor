library verilog;
use verilog.vl_types.all;
entity decoder1x2_testbench is
end decoder1x2_testbench;
