library verilog;
use verilog.vl_types.all;
entity adderC64_testbench is
end adderC64_testbench;
