../../src/verilog/signExtend12.sv