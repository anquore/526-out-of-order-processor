../../src/verilog/signExtend19.sv