../../src/verilog/mux32x64.sv