library verilog;
use verilog.vl_types.all;
entity decoder4x16_testbench is
end decoder4x16_testbench;
