../../src/verilog/decoder5x32.sv