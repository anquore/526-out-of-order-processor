../../src/verilog/D_FF.sv