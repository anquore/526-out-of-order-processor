../../src/verilog/mux_2x1_X65.sv