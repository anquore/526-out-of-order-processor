../../src/verilog/decodeStage.sv