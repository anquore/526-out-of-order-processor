library verilog;
use verilog.vl_types.all;
entity norifier_testbench is
end norifier_testbench;
