../../src/verilog/regfile.sv