../../src/verilog/NAND_MUX_2x1.sv