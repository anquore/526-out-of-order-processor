../../src/verilog/mux2_1.sv