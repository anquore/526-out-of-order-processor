../../src/verilog/commitStage.sv