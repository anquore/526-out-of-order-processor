../../src/verilog/bitSlice.sv