library verilog;
use verilog.vl_types.all;
entity signExtend19_testbench is
end signExtend19_testbench;
