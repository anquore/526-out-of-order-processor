../../src/verilog/adder64.sv