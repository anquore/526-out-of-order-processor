library verilog;
use verilog.vl_types.all;
entity multiplier_testbench is
end multiplier_testbench;
