../../src/verilog/ROB.sv