../../src/verilog/fullAdderArray63.sv