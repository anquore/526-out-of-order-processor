module registerX64(out, in, rst, clk);
	output [63:0] out;
	input [63:0] in;
	input rst, clk;
	
		D_FF r7(.q(out[7]), .d(in[7]), .reset(rst), .clk);
	D_FF r6(.q(out[6]), .d(in[6]), .reset(rst), .clk);
	D_FF r5(.q(out[5]), .d(in[5]), .reset(rst), .clk);
	D_FF r4(.q(out[4]), .d(in[4]), .reset(rst), .clk);
	D_FF r3(.q(out[3]), .d(in[3]), .reset(rst), .clk);
	D_FF r2(.q(out[2]), .d(in[2]), .reset(rst), .clk);
	D_FF r1(.q(out[1]), .d(in[1]), .reset(rst), .clk);
	D_FF r0(.q(out[0]), .d(in[0]), .reset(rst), .clk);
		D_FF r15(.q(out[15]), .d(in[15]), .reset(rst), .clk);
	D_FF r14(.q(out[14]), .d(in[14]), .reset(rst), .clk);
	D_FF r13(.q(out[13]), .d(in[13]), .reset(rst), .clk);
	D_FF r12(.q(out[12]), .d(in[12]), .reset(rst), .clk);
	D_FF r11(.q(out[11]), .d(in[11]), .reset(rst), .clk);
	D_FF r10(.q(out[10]), .d(in[10]), .reset(rst), .clk);
	D_FF r9(.q(out[9]), .d(in[9]), .reset(rst), .clk);
	D_FF r8(.q(out[8]), .d(in[8]), .reset(rst), .clk);
		D_FF r23(.q(out[23]), .d(in[23]), .reset(rst), .clk);
	D_FF r22(.q(out[22]), .d(in[22]), .reset(rst), .clk);
	D_FF r21(.q(out[21]), .d(in[21]), .reset(rst), .clk);
	D_FF r20(.q(out[20]), .d(in[20]), .reset(rst), .clk);
	D_FF r19(.q(out[19]), .d(in[19]), .reset(rst), .clk);
	D_FF r18(.q(out[18]), .d(in[18]), .reset(rst), .clk);
	D_FF r17(.q(out[17]), .d(in[17]), .reset(rst), .clk);
	D_FF r16(.q(out[16]), .d(in[16]), .reset(rst), .clk);
		D_FF r31(.q(out[31]), .d(in[31]), .reset(rst), .clk);
	D_FF r30(.q(out[30]), .d(in[30]), .reset(rst), .clk);
	D_FF r29(.q(out[29]), .d(in[29]), .reset(rst), .clk);
	D_FF r28(.q(out[28]), .d(in[28]), .reset(rst), .clk);
	D_FF r27(.q(out[27]), .d(in[27]), .reset(rst), .clk);
	D_FF r26(.q(out[26]), .d(in[26]), .reset(rst), .clk);
	D_FF r25(.q(out[25]), .d(in[25]), .reset(rst), .clk);
	D_FF r24(.q(out[24]), .d(in[24]), .reset(rst), .clk);
		D_FF r39(.q(out[39]), .d(in[39]), .reset(rst), .clk);
	D_FF r38(.q(out[38]), .d(in[38]), .reset(rst), .clk);
	D_FF r37(.q(out[37]), .d(in[37]), .reset(rst), .clk);
	D_FF r36(.q(out[36]), .d(in[36]), .reset(rst), .clk);
	D_FF r35(.q(out[35]), .d(in[35]), .reset(rst), .clk);
	D_FF r34(.q(out[34]), .d(in[34]), .reset(rst), .clk);
	D_FF r33(.q(out[33]), .d(in[33]), .reset(rst), .clk);
	D_FF r32(.q(out[32]), .d(in[32]), .reset(rst), .clk);
		D_FF r47(.q(out[47]), .d(in[47]), .reset(rst), .clk);
	D_FF r46(.q(out[46]), .d(in[46]), .reset(rst), .clk);
	D_FF r45(.q(out[45]), .d(in[45]), .reset(rst), .clk);
	D_FF r44(.q(out[44]), .d(in[44]), .reset(rst), .clk);
	D_FF r43(.q(out[43]), .d(in[43]), .reset(rst), .clk);
	D_FF r42(.q(out[42]), .d(in[42]), .reset(rst), .clk);
	D_FF r41(.q(out[41]), .d(in[41]), .reset(rst), .clk);
	D_FF r40(.q(out[40]), .d(in[40]), .reset(rst), .clk);
		D_FF r55(.q(out[55]), .d(in[55]), .reset(rst), .clk);
	D_FF r54(.q(out[54]), .d(in[54]), .reset(rst), .clk);
	D_FF r53(.q(out[53]), .d(in[53]), .reset(rst), .clk);
	D_FF r52(.q(out[52]), .d(in[52]), .reset(rst), .clk);
	D_FF r51(.q(out[51]), .d(in[51]), .reset(rst), .clk);
	D_FF r50(.q(out[50]), .d(in[50]), .reset(rst), .clk);
	D_FF r49(.q(out[49]), .d(in[49]), .reset(rst), .clk);
	D_FF r48(.q(out[48]), .d(in[48]), .reset(rst), .clk);
		D_FF r63(.q(out[63]), .d(in[63]), .reset(rst), .clk);
	D_FF r62(.q(out[62]), .d(in[62]), .reset(rst), .clk);
	D_FF r61(.q(out[61]), .d(in[61]), .reset(rst), .clk);
	D_FF r60(.q(out[60]), .d(in[60]), .reset(rst), .clk);
	D_FF r59(.q(out[59]), .d(in[59]), .reset(rst), .clk);
	D_FF r58(.q(out[58]), .d(in[58]), .reset(rst), .clk);
	D_FF r57(.q(out[57]), .d(in[57]), .reset(rst), .clk);
	D_FF r56(.q(out[56]), .d(in[56]), .reset(rst), .clk);
endmodule
