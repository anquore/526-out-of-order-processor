../../src/verilog/mux32xY.sv