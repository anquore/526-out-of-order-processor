../../src/verilog/shifter.sv