../../src/verilog/enableD_FF.sv