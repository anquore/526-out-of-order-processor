../../src/verilog/completionStage.sv