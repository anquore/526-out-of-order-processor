library verilog;
use verilog.vl_types.all;
entity shiftLeft2_testbench is
end shiftLeft2_testbench;
