../../src/verilog/headTailROB.sv