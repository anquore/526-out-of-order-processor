library verilog;
use verilog.vl_types.all;
entity mux2x64_testbench is
end mux2x64_testbench;
