../../src/verilog/mux_4x1_X64.sv