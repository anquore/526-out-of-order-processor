../../src/verilog/registerX65.sv