../../src/verilog/xnorifier.sv