library verilog;
use verilog.vl_types.all;
entity signExtend9_testbench is
end signExtend9_testbench;
