
module ROBregs ( clk_i, resets_i, decodeReadAddr1_i, decodeReadAddr2_i, 
        decodeWriteAddr_i, decodeWriteEn_i, decodeReadData1_o, 
        decodeReadData2_o, decodeWriteData_i, completionWriteAddr_i, 
        completionWriteEn_i, completionWriteData_i, commitReadAddr_i, 
        commitReadData_o );
  input [7:0] resets_i;
  input [2:0] decodeReadAddr1_i;
  input [2:0] decodeReadAddr2_i;
  input [2:0] decodeWriteAddr_i;
  output [69:0] decodeReadData1_o;
  output [69:0] decodeReadData2_o;
  input [8:0] decodeWriteData_i;
  input [2:0] completionWriteAddr_i;
  input [69:0] completionWriteData_i;
  input [2:0] commitReadAddr_i;
  output [78:0] commitReadData_o;
  input clk_i, decodeWriteEn_i, completionWriteEn_i;
  wire   n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         \managementDataOut[7][8] , \managementDataOut[7][7] ,
         \managementDataOut[7][6] , \managementDataOut[7][5] ,
         \managementDataOut[7][4] , \managementDataOut[7][3] ,
         \managementDataOut[7][2] , \managementDataOut[7][1] ,
         \managementDataOut[7][0] , \managementDataOut[6][8] ,
         \managementDataOut[6][7] , \managementDataOut[6][6] ,
         \managementDataOut[6][5] , \managementDataOut[6][4] ,
         \managementDataOut[6][3] , \managementDataOut[6][2] ,
         \managementDataOut[6][1] , \managementDataOut[6][0] ,
         \managementDataOut[5][8] , \managementDataOut[5][7] ,
         \managementDataOut[5][6] , \managementDataOut[5][5] ,
         \managementDataOut[5][4] , \managementDataOut[5][3] ,
         \managementDataOut[5][2] , \managementDataOut[5][1] ,
         \managementDataOut[5][0] , \managementDataOut[4][8] ,
         \managementDataOut[4][7] , \managementDataOut[4][6] ,
         \managementDataOut[4][5] , \managementDataOut[4][4] ,
         \managementDataOut[4][3] , \managementDataOut[4][2] ,
         \managementDataOut[4][1] , \managementDataOut[4][0] ,
         \managementDataOut[3][8] , \managementDataOut[3][7] ,
         \managementDataOut[3][6] , \managementDataOut[3][5] ,
         \managementDataOut[3][4] , \managementDataOut[3][3] ,
         \managementDataOut[3][2] , \managementDataOut[3][1] ,
         \managementDataOut[3][0] , \managementDataOut[2][8] ,
         \managementDataOut[2][7] , \managementDataOut[2][6] ,
         \managementDataOut[2][5] , \managementDataOut[2][4] ,
         \managementDataOut[2][3] , \managementDataOut[2][2] ,
         \managementDataOut[2][1] , \managementDataOut[2][0] ,
         \managementDataOut[1][8] , \managementDataOut[1][7] ,
         \managementDataOut[1][6] , \managementDataOut[1][5] ,
         \managementDataOut[1][4] , \managementDataOut[1][3] ,
         \managementDataOut[1][2] , \managementDataOut[1][1] ,
         \managementDataOut[1][0] , \managementDataOut[0][8] ,
         \managementDataOut[0][7] , \managementDataOut[0][6] ,
         \managementDataOut[0][5] , \managementDataOut[0][4] ,
         \managementDataOut[0][3] , \managementDataOut[0][2] ,
         \managementDataOut[0][1] , \managementDataOut[0][0] ,
         \completionDataOut[7][69] , \completionDataOut[7][68] ,
         \completionDataOut[7][67] , \completionDataOut[7][66] ,
         \completionDataOut[7][65] , \completionDataOut[7][64] ,
         \completionDataOut[7][63] , \completionDataOut[7][62] ,
         \completionDataOut[7][61] , \completionDataOut[7][60] ,
         \completionDataOut[7][59] , \completionDataOut[7][58] ,
         \completionDataOut[7][57] , \completionDataOut[7][56] ,
         \completionDataOut[7][55] , \completionDataOut[7][54] ,
         \completionDataOut[7][53] , \completionDataOut[7][52] ,
         \completionDataOut[7][51] , \completionDataOut[7][50] ,
         \completionDataOut[7][49] , \completionDataOut[7][48] ,
         \completionDataOut[7][47] , \completionDataOut[7][46] ,
         \completionDataOut[7][45] , \completionDataOut[7][44] ,
         \completionDataOut[7][43] , \completionDataOut[7][42] ,
         \completionDataOut[7][41] , \completionDataOut[7][40] ,
         \completionDataOut[7][39] , \completionDataOut[7][38] ,
         \completionDataOut[7][37] , \completionDataOut[7][36] ,
         \completionDataOut[7][35] , \completionDataOut[7][34] ,
         \completionDataOut[7][33] , \completionDataOut[7][32] ,
         \completionDataOut[7][31] , \completionDataOut[7][30] ,
         \completionDataOut[7][29] , \completionDataOut[7][28] ,
         \completionDataOut[7][27] , \completionDataOut[7][26] ,
         \completionDataOut[7][25] , \completionDataOut[7][24] ,
         \completionDataOut[7][23] , \completionDataOut[7][22] ,
         \completionDataOut[7][21] , \completionDataOut[7][20] ,
         \completionDataOut[7][19] , \completionDataOut[7][18] ,
         \completionDataOut[7][17] , \completionDataOut[7][16] ,
         \completionDataOut[7][15] , \completionDataOut[7][14] ,
         \completionDataOut[7][13] , \completionDataOut[7][12] ,
         \completionDataOut[7][11] , \completionDataOut[7][10] ,
         \completionDataOut[7][9] , \completionDataOut[7][8] ,
         \completionDataOut[7][7] , \completionDataOut[7][6] ,
         \completionDataOut[7][5] , \completionDataOut[7][4] ,
         \completionDataOut[7][3] , \completionDataOut[7][2] ,
         \completionDataOut[7][1] , \completionDataOut[7][0] ,
         \completionDataOut[6][69] , \completionDataOut[6][68] ,
         \completionDataOut[6][67] , \completionDataOut[6][66] ,
         \completionDataOut[6][65] , \completionDataOut[6][64] ,
         \completionDataOut[6][63] , \completionDataOut[6][62] ,
         \completionDataOut[6][61] , \completionDataOut[6][60] ,
         \completionDataOut[6][59] , \completionDataOut[6][58] ,
         \completionDataOut[6][57] , \completionDataOut[6][56] ,
         \completionDataOut[6][55] , \completionDataOut[6][54] ,
         \completionDataOut[6][53] , \completionDataOut[6][52] ,
         \completionDataOut[6][51] , \completionDataOut[6][50] ,
         \completionDataOut[6][49] , \completionDataOut[6][48] ,
         \completionDataOut[6][47] , \completionDataOut[6][46] ,
         \completionDataOut[6][45] , \completionDataOut[6][44] ,
         \completionDataOut[6][43] , \completionDataOut[6][42] ,
         \completionDataOut[6][41] , \completionDataOut[6][40] ,
         \completionDataOut[6][39] , \completionDataOut[6][38] ,
         \completionDataOut[6][37] , \completionDataOut[6][36] ,
         \completionDataOut[6][35] , \completionDataOut[6][34] ,
         \completionDataOut[6][33] , \completionDataOut[6][32] ,
         \completionDataOut[6][31] , \completionDataOut[6][30] ,
         \completionDataOut[6][29] , \completionDataOut[6][28] ,
         \completionDataOut[6][27] , \completionDataOut[6][26] ,
         \completionDataOut[6][25] , \completionDataOut[6][24] ,
         \completionDataOut[6][23] , \completionDataOut[6][22] ,
         \completionDataOut[6][21] , \completionDataOut[6][20] ,
         \completionDataOut[6][19] , \completionDataOut[6][18] ,
         \completionDataOut[6][17] , \completionDataOut[6][16] ,
         \completionDataOut[6][15] , \completionDataOut[6][14] ,
         \completionDataOut[6][13] , \completionDataOut[6][12] ,
         \completionDataOut[6][11] , \completionDataOut[6][10] ,
         \completionDataOut[6][9] , \completionDataOut[6][8] ,
         \completionDataOut[6][7] , \completionDataOut[6][6] ,
         \completionDataOut[6][5] , \completionDataOut[6][4] ,
         \completionDataOut[6][3] , \completionDataOut[6][2] ,
         \completionDataOut[6][1] , \completionDataOut[6][0] ,
         \completionDataOut[5][69] , \completionDataOut[5][68] ,
         \completionDataOut[5][67] , \completionDataOut[5][66] ,
         \completionDataOut[5][65] , \completionDataOut[5][64] ,
         \completionDataOut[5][63] , \completionDataOut[5][62] ,
         \completionDataOut[5][61] , \completionDataOut[5][60] ,
         \completionDataOut[5][59] , \completionDataOut[5][58] ,
         \completionDataOut[5][57] , \completionDataOut[5][56] ,
         \completionDataOut[5][55] , \completionDataOut[5][54] ,
         \completionDataOut[5][53] , \completionDataOut[5][52] ,
         \completionDataOut[5][51] , \completionDataOut[5][50] ,
         \completionDataOut[5][49] , \completionDataOut[5][48] ,
         \completionDataOut[5][47] , \completionDataOut[5][46] ,
         \completionDataOut[5][45] , \completionDataOut[5][44] ,
         \completionDataOut[5][43] , \completionDataOut[5][42] ,
         \completionDataOut[5][41] , \completionDataOut[5][40] ,
         \completionDataOut[5][39] , \completionDataOut[5][38] ,
         \completionDataOut[5][37] , \completionDataOut[5][36] ,
         \completionDataOut[5][35] , \completionDataOut[5][34] ,
         \completionDataOut[5][33] , \completionDataOut[5][32] ,
         \completionDataOut[5][31] , \completionDataOut[5][30] ,
         \completionDataOut[5][29] , \completionDataOut[5][28] ,
         \completionDataOut[5][27] , \completionDataOut[5][26] ,
         \completionDataOut[5][25] , \completionDataOut[5][24] ,
         \completionDataOut[5][23] , \completionDataOut[5][22] ,
         \completionDataOut[5][21] , \completionDataOut[5][20] ,
         \completionDataOut[5][19] , \completionDataOut[5][18] ,
         \completionDataOut[5][17] , \completionDataOut[5][16] ,
         \completionDataOut[5][15] , \completionDataOut[5][14] ,
         \completionDataOut[5][13] , \completionDataOut[5][12] ,
         \completionDataOut[5][11] , \completionDataOut[5][10] ,
         \completionDataOut[5][9] , \completionDataOut[5][8] ,
         \completionDataOut[5][7] , \completionDataOut[5][6] ,
         \completionDataOut[5][5] , \completionDataOut[5][4] ,
         \completionDataOut[5][3] , \completionDataOut[5][2] ,
         \completionDataOut[5][1] , \completionDataOut[5][0] ,
         \completionDataOut[4][69] , \completionDataOut[4][68] ,
         \completionDataOut[4][67] , \completionDataOut[4][66] ,
         \completionDataOut[4][65] , \completionDataOut[4][64] ,
         \completionDataOut[4][63] , \completionDataOut[4][62] ,
         \completionDataOut[4][61] , \completionDataOut[4][60] ,
         \completionDataOut[4][59] , \completionDataOut[4][58] ,
         \completionDataOut[4][57] , \completionDataOut[4][56] ,
         \completionDataOut[4][55] , \completionDataOut[4][54] ,
         \completionDataOut[4][53] , \completionDataOut[4][52] ,
         \completionDataOut[4][51] , \completionDataOut[4][50] ,
         \completionDataOut[4][49] , \completionDataOut[4][48] ,
         \completionDataOut[4][47] , \completionDataOut[4][46] ,
         \completionDataOut[4][45] , \completionDataOut[4][44] ,
         \completionDataOut[4][43] , \completionDataOut[4][42] ,
         \completionDataOut[4][41] , \completionDataOut[4][40] ,
         \completionDataOut[4][39] , \completionDataOut[4][38] ,
         \completionDataOut[4][37] , \completionDataOut[4][36] ,
         \completionDataOut[4][35] , \completionDataOut[4][34] ,
         \completionDataOut[4][33] , \completionDataOut[4][32] ,
         \completionDataOut[4][31] , \completionDataOut[4][30] ,
         \completionDataOut[4][29] , \completionDataOut[4][28] ,
         \completionDataOut[4][27] , \completionDataOut[4][26] ,
         \completionDataOut[4][25] , \completionDataOut[4][24] ,
         \completionDataOut[4][23] , \completionDataOut[4][22] ,
         \completionDataOut[4][21] , \completionDataOut[4][20] ,
         \completionDataOut[4][19] , \completionDataOut[4][18] ,
         \completionDataOut[4][17] , \completionDataOut[4][16] ,
         \completionDataOut[4][15] , \completionDataOut[4][14] ,
         \completionDataOut[4][13] , \completionDataOut[4][12] ,
         \completionDataOut[4][11] , \completionDataOut[4][10] ,
         \completionDataOut[4][9] , \completionDataOut[4][8] ,
         \completionDataOut[4][7] , \completionDataOut[4][6] ,
         \completionDataOut[4][5] , \completionDataOut[4][4] ,
         \completionDataOut[4][3] , \completionDataOut[4][2] ,
         \completionDataOut[4][1] , \completionDataOut[4][0] ,
         \completionDataOut[3][69] , \completionDataOut[3][68] ,
         \completionDataOut[3][67] , \completionDataOut[3][66] ,
         \completionDataOut[3][65] , \completionDataOut[3][64] ,
         \completionDataOut[3][63] , \completionDataOut[3][62] ,
         \completionDataOut[3][61] , \completionDataOut[3][60] ,
         \completionDataOut[3][59] , \completionDataOut[3][58] ,
         \completionDataOut[3][57] , \completionDataOut[3][56] ,
         \completionDataOut[3][55] , \completionDataOut[3][54] ,
         \completionDataOut[3][53] , \completionDataOut[3][52] ,
         \completionDataOut[3][51] , \completionDataOut[3][50] ,
         \completionDataOut[3][49] , \completionDataOut[3][48] ,
         \completionDataOut[3][47] , \completionDataOut[3][46] ,
         \completionDataOut[3][45] , \completionDataOut[3][44] ,
         \completionDataOut[3][43] , \completionDataOut[3][42] ,
         \completionDataOut[3][41] , \completionDataOut[3][40] ,
         \completionDataOut[3][39] , \completionDataOut[3][38] ,
         \completionDataOut[3][37] , \completionDataOut[3][36] ,
         \completionDataOut[3][35] , \completionDataOut[3][34] ,
         \completionDataOut[3][33] , \completionDataOut[3][32] ,
         \completionDataOut[3][31] , \completionDataOut[3][30] ,
         \completionDataOut[3][29] , \completionDataOut[3][28] ,
         \completionDataOut[3][27] , \completionDataOut[3][26] ,
         \completionDataOut[3][25] , \completionDataOut[3][24] ,
         \completionDataOut[3][23] , \completionDataOut[3][22] ,
         \completionDataOut[3][21] , \completionDataOut[3][20] ,
         \completionDataOut[3][19] , \completionDataOut[3][18] ,
         \completionDataOut[3][17] , \completionDataOut[3][16] ,
         \completionDataOut[3][15] , \completionDataOut[3][14] ,
         \completionDataOut[3][13] , \completionDataOut[3][12] ,
         \completionDataOut[3][11] , \completionDataOut[3][10] ,
         \completionDataOut[3][9] , \completionDataOut[3][8] ,
         \completionDataOut[3][7] , \completionDataOut[3][6] ,
         \completionDataOut[3][5] , \completionDataOut[3][4] ,
         \completionDataOut[3][3] , \completionDataOut[3][2] ,
         \completionDataOut[3][1] , \completionDataOut[3][0] ,
         \completionDataOut[2][69] , \completionDataOut[2][68] ,
         \completionDataOut[2][67] , \completionDataOut[2][66] ,
         \completionDataOut[2][65] , \completionDataOut[2][64] ,
         \completionDataOut[2][63] , \completionDataOut[2][62] ,
         \completionDataOut[2][61] , \completionDataOut[2][60] ,
         \completionDataOut[2][59] , \completionDataOut[2][58] ,
         \completionDataOut[2][57] , \completionDataOut[2][56] ,
         \completionDataOut[2][55] , \completionDataOut[2][54] ,
         \completionDataOut[2][53] , \completionDataOut[2][52] ,
         \completionDataOut[2][51] , \completionDataOut[2][50] ,
         \completionDataOut[2][49] , \completionDataOut[2][48] ,
         \completionDataOut[2][47] , \completionDataOut[2][46] ,
         \completionDataOut[2][45] , \completionDataOut[2][44] ,
         \completionDataOut[2][43] , \completionDataOut[2][42] ,
         \completionDataOut[2][41] , \completionDataOut[2][40] ,
         \completionDataOut[2][39] , \completionDataOut[2][38] ,
         \completionDataOut[2][37] , \completionDataOut[2][36] ,
         \completionDataOut[2][35] , \completionDataOut[2][34] ,
         \completionDataOut[2][33] , \completionDataOut[2][32] ,
         \completionDataOut[2][31] , \completionDataOut[2][30] ,
         \completionDataOut[2][29] , \completionDataOut[2][28] ,
         \completionDataOut[2][27] , \completionDataOut[2][26] ,
         \completionDataOut[2][25] , \completionDataOut[2][24] ,
         \completionDataOut[2][23] , \completionDataOut[2][22] ,
         \completionDataOut[2][21] , \completionDataOut[2][20] ,
         \completionDataOut[2][19] , \completionDataOut[2][18] ,
         \completionDataOut[2][17] , \completionDataOut[2][16] ,
         \completionDataOut[2][15] , \completionDataOut[2][14] ,
         \completionDataOut[2][13] , \completionDataOut[2][12] ,
         \completionDataOut[2][11] , \completionDataOut[2][10] ,
         \completionDataOut[2][9] , \completionDataOut[2][8] ,
         \completionDataOut[2][7] , \completionDataOut[2][6] ,
         \completionDataOut[2][5] , \completionDataOut[2][4] ,
         \completionDataOut[2][3] , \completionDataOut[2][2] ,
         \completionDataOut[2][1] , \completionDataOut[2][0] ,
         \completionDataOut[1][69] , \completionDataOut[1][68] ,
         \completionDataOut[1][67] , \completionDataOut[1][66] ,
         \completionDataOut[1][65] , \completionDataOut[1][64] ,
         \completionDataOut[1][63] , \completionDataOut[1][62] ,
         \completionDataOut[1][61] , \completionDataOut[1][60] ,
         \completionDataOut[1][59] , \completionDataOut[1][58] ,
         \completionDataOut[1][57] , \completionDataOut[1][56] ,
         \completionDataOut[1][55] , \completionDataOut[1][54] ,
         \completionDataOut[1][53] , \completionDataOut[1][52] ,
         \completionDataOut[1][51] , \completionDataOut[1][50] ,
         \completionDataOut[1][49] , \completionDataOut[1][48] ,
         \completionDataOut[1][47] , \completionDataOut[1][46] ,
         \completionDataOut[1][45] , \completionDataOut[1][44] ,
         \completionDataOut[1][43] , \completionDataOut[1][42] ,
         \completionDataOut[1][41] , \completionDataOut[1][40] ,
         \completionDataOut[1][39] , \completionDataOut[1][38] ,
         \completionDataOut[1][37] , \completionDataOut[1][36] ,
         \completionDataOut[1][35] , \completionDataOut[1][34] ,
         \completionDataOut[1][33] , \completionDataOut[1][32] ,
         \completionDataOut[1][31] , \completionDataOut[1][30] ,
         \completionDataOut[1][29] , \completionDataOut[1][28] ,
         \completionDataOut[1][27] , \completionDataOut[1][26] ,
         \completionDataOut[1][25] , \completionDataOut[1][24] ,
         \completionDataOut[1][23] , \completionDataOut[1][22] ,
         \completionDataOut[1][21] , \completionDataOut[1][20] ,
         \completionDataOut[1][19] , \completionDataOut[1][18] ,
         \completionDataOut[1][17] , \completionDataOut[1][16] ,
         \completionDataOut[1][15] , \completionDataOut[1][14] ,
         \completionDataOut[1][13] , \completionDataOut[1][12] ,
         \completionDataOut[1][11] , \completionDataOut[1][10] ,
         \completionDataOut[1][9] , \completionDataOut[1][8] ,
         \completionDataOut[1][7] , \completionDataOut[1][6] ,
         \completionDataOut[1][5] , \completionDataOut[1][4] ,
         \completionDataOut[1][3] , \completionDataOut[1][2] ,
         \completionDataOut[1][1] , \completionDataOut[1][0] ,
         \completionDataOut[0][69] , \completionDataOut[0][68] ,
         \completionDataOut[0][67] , \completionDataOut[0][66] ,
         \completionDataOut[0][65] , \completionDataOut[0][64] ,
         \completionDataOut[0][63] , \completionDataOut[0][62] ,
         \completionDataOut[0][61] , \completionDataOut[0][60] ,
         \completionDataOut[0][59] , \completionDataOut[0][58] ,
         \completionDataOut[0][57] , \completionDataOut[0][56] ,
         \completionDataOut[0][55] , \completionDataOut[0][54] ,
         \completionDataOut[0][53] , \completionDataOut[0][52] ,
         \completionDataOut[0][51] , \completionDataOut[0][50] ,
         \completionDataOut[0][49] , \completionDataOut[0][48] ,
         \completionDataOut[0][47] , \completionDataOut[0][46] ,
         \completionDataOut[0][45] , \completionDataOut[0][44] ,
         \completionDataOut[0][43] , \completionDataOut[0][42] ,
         \completionDataOut[0][41] , \completionDataOut[0][40] ,
         \completionDataOut[0][39] , \completionDataOut[0][38] ,
         \completionDataOut[0][37] , \completionDataOut[0][36] ,
         \completionDataOut[0][35] , \completionDataOut[0][34] ,
         \completionDataOut[0][33] , \completionDataOut[0][32] ,
         \completionDataOut[0][31] , \completionDataOut[0][30] ,
         \completionDataOut[0][29] , \completionDataOut[0][28] ,
         \completionDataOut[0][27] , \completionDataOut[0][26] ,
         \completionDataOut[0][25] , \completionDataOut[0][24] ,
         \completionDataOut[0][23] , \completionDataOut[0][22] ,
         \completionDataOut[0][21] , \completionDataOut[0][20] ,
         \completionDataOut[0][19] , \completionDataOut[0][18] ,
         \completionDataOut[0][17] , \completionDataOut[0][16] ,
         \completionDataOut[0][15] , \completionDataOut[0][14] ,
         \completionDataOut[0][13] , \completionDataOut[0][12] ,
         \completionDataOut[0][11] , \completionDataOut[0][10] ,
         \completionDataOut[0][9] , \completionDataOut[0][8] ,
         \completionDataOut[0][7] , \completionDataOut[0][6] ,
         \completionDataOut[0][5] , \completionDataOut[0][4] ,
         \completionDataOut[0][3] , \completionDataOut[0][2] ,
         \completionDataOut[0][1] , \completionDataOut[0][0] ,
         \eachManagementReg[2].managementReg/eachEnDff[0].enDff/theFlop/N3 ,
         \eachManagementReg[2].managementReg/eachEnDff[1].enDff/theFlop/N3 ,
         \eachManagementReg[2].managementReg/eachEnDff[2].enDff/theFlop/N3 ,
         \eachManagementReg[2].managementReg/eachEnDff[3].enDff/theFlop/N3 ,
         \eachManagementReg[2].managementReg/eachEnDff[4].enDff/theFlop/N3 ,
         \eachManagementReg[2].managementReg/eachEnDff[5].enDff/theFlop/N3 ,
         \eachManagementReg[2].managementReg/eachEnDff[6].enDff/theFlop/N3 ,
         \eachManagementReg[2].managementReg/eachEnDff[7].enDff/theFlop/N3 ,
         \eachManagementReg[2].managementReg/eachEnDff[8].enDff/theFlop/N3 ,
         \eachManagementReg[3].managementReg/eachEnDff[0].enDff/theFlop/N3 ,
         \eachManagementReg[3].managementReg/eachEnDff[1].enDff/theFlop/N3 ,
         \eachManagementReg[3].managementReg/eachEnDff[2].enDff/theFlop/N3 ,
         \eachManagementReg[3].managementReg/eachEnDff[3].enDff/theFlop/N3 ,
         \eachManagementReg[3].managementReg/eachEnDff[4].enDff/theFlop/N3 ,
         \eachManagementReg[3].managementReg/eachEnDff[5].enDff/theFlop/N3 ,
         \eachManagementReg[3].managementReg/eachEnDff[6].enDff/theFlop/N3 ,
         \eachManagementReg[3].managementReg/eachEnDff[7].enDff/theFlop/N3 ,
         \eachManagementReg[3].managementReg/eachEnDff[8].enDff/theFlop/N3 ,
         \eachManagementReg[5].managementReg/eachEnDff[0].enDff/theFlop/N3 ,
         \eachManagementReg[5].managementReg/eachEnDff[1].enDff/theFlop/N3 ,
         \eachManagementReg[5].managementReg/eachEnDff[2].enDff/theFlop/N3 ,
         \eachManagementReg[5].managementReg/eachEnDff[3].enDff/theFlop/N3 ,
         \eachManagementReg[5].managementReg/eachEnDff[4].enDff/theFlop/N3 ,
         \eachManagementReg[5].managementReg/eachEnDff[5].enDff/theFlop/N3 ,
         \eachManagementReg[5].managementReg/eachEnDff[6].enDff/theFlop/N3 ,
         \eachManagementReg[5].managementReg/eachEnDff[7].enDff/theFlop/N3 ,
         \eachManagementReg[5].managementReg/eachEnDff[8].enDff/theFlop/N3 ,
         \eachManagementReg[6].managementReg/eachEnDff[0].enDff/theFlop/N3 ,
         \eachManagementReg[6].managementReg/eachEnDff[1].enDff/theFlop/N3 ,
         \eachManagementReg[6].managementReg/eachEnDff[2].enDff/theFlop/N3 ,
         \eachManagementReg[6].managementReg/eachEnDff[3].enDff/theFlop/N3 ,
         \eachManagementReg[6].managementReg/eachEnDff[4].enDff/theFlop/N3 ,
         \eachManagementReg[6].managementReg/eachEnDff[5].enDff/theFlop/N3 ,
         \eachManagementReg[6].managementReg/eachEnDff[6].enDff/theFlop/N3 ,
         \eachManagementReg[6].managementReg/eachEnDff[7].enDff/theFlop/N3 ,
         \eachManagementReg[6].managementReg/eachEnDff[8].enDff/theFlop/N3 ,
         \eachManagementReg[7].managementReg/eachEnDff[0].enDff/theFlop/N3 ,
         \eachManagementReg[7].managementReg/eachEnDff[1].enDff/theFlop/N3 ,
         \eachManagementReg[7].managementReg/eachEnDff[2].enDff/theFlop/N3 ,
         \eachManagementReg[7].managementReg/eachEnDff[3].enDff/theFlop/N3 ,
         \eachManagementReg[7].managementReg/eachEnDff[4].enDff/theFlop/N3 ,
         \eachManagementReg[7].managementReg/eachEnDff[5].enDff/theFlop/N3 ,
         \eachManagementReg[7].managementReg/eachEnDff[6].enDff/theFlop/N3 ,
         \eachManagementReg[7].managementReg/eachEnDff[7].enDff/theFlop/N3 ,
         \eachManagementReg[7].managementReg/eachEnDff[8].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[0].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[1].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[2].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[3].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[4].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[5].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[6].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[7].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[8].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[9].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[10].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[11].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[12].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[13].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[14].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[15].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[16].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[17].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[18].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[19].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[20].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[21].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[22].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[23].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[24].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[25].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[26].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[27].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[28].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[29].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[30].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[31].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[32].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[33].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[34].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[35].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[36].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[37].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[38].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[39].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[40].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[41].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[42].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[43].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[44].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[45].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[46].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[47].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[48].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[49].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[50].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[51].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[52].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[53].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[54].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[55].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[56].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[57].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[58].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[59].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[60].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[61].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[62].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[63].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[64].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[65].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[66].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[67].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[68].enDff/theFlop/N3 ,
         \eachCompletionReg[2].completionReg/eachEnDff[69].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[0].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[1].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[2].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[3].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[4].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[5].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[6].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[7].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[8].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[9].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[10].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[11].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[12].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[13].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[14].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[15].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[16].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[17].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[18].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[19].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[20].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[21].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[22].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[23].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[24].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[25].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[26].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[27].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[28].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[29].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[30].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[31].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[32].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[33].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[34].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[35].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[36].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[37].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[38].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[39].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[40].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[41].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[42].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[43].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[44].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[45].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[46].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[47].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[48].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[49].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[50].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[51].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[52].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[53].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[54].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[55].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[56].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[57].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[58].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[59].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[60].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[61].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[62].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[63].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[64].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[65].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[66].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[67].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[68].enDff/theFlop/N3 ,
         \eachCompletionReg[3].completionReg/eachEnDff[69].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[0].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[1].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[2].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[3].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[4].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[5].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[6].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[7].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[8].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[9].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[10].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[11].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[12].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[13].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[14].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[15].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[16].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[17].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[18].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[19].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[20].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[21].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[22].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[23].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[24].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[25].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[26].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[27].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[28].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[29].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[30].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[31].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[32].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[33].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[34].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[35].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[36].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[37].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[38].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[39].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[40].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[41].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[42].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[43].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[44].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[45].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[46].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[47].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[48].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[49].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[50].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[51].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[52].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[53].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[54].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[55].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[56].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[57].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[58].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[59].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[60].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[61].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[62].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[63].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[64].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[65].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[66].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[67].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[68].enDff/theFlop/N3 ,
         \eachCompletionReg[5].completionReg/eachEnDff[69].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[0].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[1].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[2].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[3].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[4].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[5].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[6].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[7].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[8].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[9].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[10].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[11].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[12].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[13].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[14].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[15].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[16].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[17].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[18].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[19].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[20].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[21].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[22].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[23].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[24].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[25].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[26].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[27].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[28].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[29].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[30].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[31].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[32].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[33].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[34].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[35].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[36].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[37].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[38].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[39].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[40].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[41].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[42].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[43].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[44].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[45].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[46].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[47].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[48].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[49].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[50].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[51].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[52].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[53].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[54].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[55].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[56].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[57].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[58].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[59].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[60].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[61].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[62].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[63].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[64].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[65].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[66].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[67].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[68].enDff/theFlop/N3 ,
         \eachCompletionReg[6].completionReg/eachEnDff[69].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[0].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[1].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[2].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[3].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[4].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[5].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[6].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[7].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[8].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[9].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[10].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[11].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[12].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[13].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[14].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[15].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[16].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[17].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[18].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[19].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[20].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[21].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[22].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[23].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[24].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[25].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[26].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[27].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[28].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[29].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[30].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[31].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[32].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[33].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[34].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[35].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[36].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[37].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[38].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[39].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[40].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[41].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[42].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[43].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[44].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[45].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[46].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[47].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[48].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[49].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[50].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[51].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[52].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[53].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[54].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[55].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[56].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[57].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[58].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[59].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[60].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[61].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[62].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[63].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[64].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[65].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[66].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[67].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[68].enDff/theFlop/N3 ,
         \eachCompletionReg[7].completionReg/eachEnDff[69].enDff/theFlop/N3 ,
         n1, n2, n3, n4, n5, n6, n7, n30, n49, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060;

  DFQD1 \eachManagementReg[3].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[3].managementReg/eachEnDff[0].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[3][0] ) );
  DFQD1 \eachManagementReg[3].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[3].managementReg/eachEnDff[1].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[3][1] ) );
  DFQD1 \eachManagementReg[3].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[3].managementReg/eachEnDff[4].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[3][4] ) );
  DFQD1 \eachManagementReg[3].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[3].managementReg/eachEnDff[5].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[3][5] ) );
  DFQD1 \eachManagementReg[3].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[3].managementReg/eachEnDff[6].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[3][6] ) );
  DFQD1 \eachManagementReg[3].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[3].managementReg/eachEnDff[8].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[3][8] ) );
  DFQD1 \eachManagementReg[5].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[5].managementReg/eachEnDff[2].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[5][2] ) );
  DFQD1 \eachManagementReg[5].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[5].managementReg/eachEnDff[3].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[5][3] ) );
  DFQD1 \eachManagementReg[5].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[5].managementReg/eachEnDff[4].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[5][4] ) );
  DFQD1 \eachManagementReg[5].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[5].managementReg/eachEnDff[5].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[5][5] ) );
  DFQD1 \eachManagementReg[5].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[5].managementReg/eachEnDff[6].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[5][6] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .CN(n1247), .D(completionWriteData_i[45]), .E(n61), .CP(clk_i), .Q(
        \completionDataOut[0][45] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .CN(n68), .D(completionWriteData_i[45]), .E(n59), .CP(clk_i), .Q(
        \completionDataOut[4][45] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .CN(n51), .D(completionWriteData_i[69]), .E(n44), .CP(clk_i), .Q(
        \completionDataOut[4][69] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .CN(n3), .D(completionWriteData_i[57]), .E(n178), .CP(clk_i), .Q(
        \completionDataOut[4][57] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .CN(n190), .D(completionWriteData_i[55]), .E(n46), .CP(clk_i), .Q(
        \completionDataOut[4][55] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .CN(n78), .D(completionWriteData_i[69]), .E(n1257), .CP(clk_i), .Q(
        \completionDataOut[1][69] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .CN(n95), .D(completionWriteData_i[69]), .E(n45), .CP(clk_i), .Q(
        \completionDataOut[0][69] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .CN(n84), .D(completionWriteData_i[57]), .E(n182), .CP(clk_i), .Q(
        \completionDataOut[0][57] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .CN(n1248), .D(completionWriteData_i[55]), .E(n47), .CP(clk_i), .Q(
        \completionDataOut[0][55] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .CN(n189), .D(completionWriteData_i[6]), .E(n58), .CP(clk_i), .Q(
        \completionDataOut[4][6] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .CN(n53), .D(completionWriteData_i[44]), .E(n60), .CP(clk_i), .Q(
        \completionDataOut[0][44] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .CN(n85), .D(completionWriteData_i[43]), .E(n181), .CP(clk_i), .Q(
        \completionDataOut[0][43] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .CN(n84), .D(completionWriteData_i[42]), .E(n90), .CP(clk_i), .Q(
        \completionDataOut[0][42] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .CN(n96), .D(completionWriteData_i[41]), .E(n184), .CP(clk_i), .Q(
        \completionDataOut[0][41] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .CN(n86), .D(completionWriteData_i[40]), .E(n75), .CP(clk_i), .Q(
        \completionDataOut[0][40] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .CN(n192), .D(completionWriteData_i[68]), .E(n60), .CP(clk_i), .Q(
        \completionDataOut[0][68] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .CN(n85), .D(completionWriteData_i[67]), .E(n76), .CP(clk_i), .Q(
        \completionDataOut[0][67] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .CN(n5), .D(completionWriteData_i[68]), .E(n1259), .CP(clk_i), .Q(
        \completionDataOut[1][68] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .CN(n92), .D(completionWriteData_i[67]), .E(n1257), .CP(clk_i), .Q(
        \completionDataOut[1][67] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .CN(n63), .D(completionWriteData_i[66]), .E(n1259), .CP(clk_i), .Q(
        \completionDataOut[1][66] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .CN(n84), .D(completionWriteData_i[48]), .E(n90), .CP(clk_i), .Q(
        \completionDataOut[0][48] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .CN(n1248), .D(completionWriteData_i[51]), .E(n184), .CP(clk_i), .Q(
        \completionDataOut[0][51] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .CN(n83), .D(completionWriteData_i[50]), .E(n183), .CP(clk_i), .Q(
        \completionDataOut[0][50] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .CN(n92), .D(completionWriteData_i[51]), .E(n1261), .CP(clk_i), .Q(
        \completionDataOut[1][51] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .CN(n50), .D(completionWriteData_i[50]), .E(n1261), .CP(clk_i), .Q(
        \completionDataOut[1][50] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .CN(n91), .D(completionWriteData_i[49]), .E(n1261), .CP(clk_i), .Q(
        \completionDataOut[1][49] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .CN(n80), .D(completionWriteData_i[48]), .E(n1261), .CP(clk_i), .Q(
        \completionDataOut[1][48] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .CN(n66), .D(completionWriteData_i[44]), .E(n177), .CP(clk_i), .Q(
        \completionDataOut[4][44] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .CN(n67), .D(completionWriteData_i[43]), .E(n88), .CP(clk_i), .Q(
        \completionDataOut[4][43] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .CN(n93), .D(completionWriteData_i[41]), .E(n180), .CP(clk_i), .Q(
        \completionDataOut[4][41] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .CN(n94), .D(completionWriteData_i[52]), .E(n73), .CP(clk_i), .Q(
        \completionDataOut[4][52] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .CN(n82), .D(completionWriteData_i[9]), .E(n58), .CP(clk_i), .Q(
        \completionDataOut[4][9] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .CN(n69), .D(completionWriteData_i[8]), .E(n74), .CP(clk_i), .Q(
        \completionDataOut[4][8] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .CN(n42), .D(completionWriteData_i[7]), .E(n88), .CP(clk_i), .Q(
        \completionDataOut[4][7] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .CN(n189), .D(completionWriteData_i[5]), .E(n180), .CP(clk_i), .Q(
        \completionDataOut[4][5] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .CN(n82), .D(completionWriteData_i[4]), .E(n179), .CP(clk_i), .Q(
        \completionDataOut[4][4] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .CN(n68), .D(completionWriteData_i[53]), .E(n180), .CP(clk_i), .Q(
        \completionDataOut[4][53] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .CN(n69), .D(completionWriteData_i[3]), .E(n87), .CP(clk_i), .Q(
        \completionDataOut[4][3] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .CN(n42), .D(completionWriteData_i[2]), .E(n179), .CP(clk_i), .Q(
        \completionDataOut[4][2] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .CN(n3), .D(completionWriteData_i[1]), .E(n88), .CP(clk_i), .Q(
        \completionDataOut[4][1] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .CN(n189), .D(completionWriteData_i[0]), .E(n46), .CP(clk_i), .Q(
        \completionDataOut[4][0] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .CN(n81), .D(completionWriteData_i[42]), .E(n87), .CP(clk_i), .Q(
        \completionDataOut[4][42] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .CN(n66), .D(completionWriteData_i[40]), .E(n88), .CP(clk_i), .Q(
        \completionDataOut[4][40] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .CN(n51), .D(completionWriteData_i[68]), .E(n178), .CP(clk_i), .Q(
        \completionDataOut[4][68] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .CN(n67), .D(completionWriteData_i[67]), .E(n180), .CP(clk_i), .Q(
        \completionDataOut[4][67] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .CN(n69), .D(completionWriteData_i[66]), .E(n87), .CP(clk_i), .Q(
        \completionDataOut[4][66] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .CN(n189), .D(completionWriteData_i[65]), .E(n74), .CP(clk_i), .Q(
        \completionDataOut[4][65] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .CN(n93), .D(completionWriteData_i[64]), .E(n59), .CP(clk_i), .Q(
        \completionDataOut[4][64] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .CN(n67), .D(completionWriteData_i[56]), .E(n179), .CP(clk_i), .Q(
        \completionDataOut[4][56] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .CN(n52), .D(completionWriteData_i[54]), .E(n44), .CP(clk_i), .Q(
        \completionDataOut[4][54] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .CN(n66), .D(completionWriteData_i[51]), .E(n179), .CP(clk_i), .Q(
        \completionDataOut[4][51] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .CN(n52), .D(completionWriteData_i[50]), .E(n59), .CP(clk_i), .Q(
        \completionDataOut[4][50] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .CN(n190), .D(completionWriteData_i[49]), .E(n179), .CP(clk_i), .Q(
        \completionDataOut[4][49] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .CN(n81), .D(completionWriteData_i[48]), .E(n73), .CP(clk_i), .Q(
        \completionDataOut[4][48] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .CN(n69), .D(completionWriteData_i[47]), .E(n177), .CP(clk_i), .Q(
        \completionDataOut[4][47] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .CN(n64), .D(completionWriteData_i[65]), .E(n1256), .CP(clk_i), .Q(
        \completionDataOut[1][65] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .CN(n68), .D(completionWriteData_i[46]), .E(n177), .CP(clk_i), .Q(
        \completionDataOut[4][46] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .CN(n186), .D(completionWriteData_i[9]), .E(n1255), .CP(clk_i), .Q(
        \completionDataOut[1][9] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .CN(n186), .D(completionWriteData_i[8]), .E(n1255), .CP(clk_i), .Q(
        \completionDataOut[1][8] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .CN(n64), .D(completionWriteData_i[7]), .E(n1255), .CP(clk_i), .Q(
        \completionDataOut[1][7] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .CN(n78), .D(completionWriteData_i[6]), .E(n1255), .CP(clk_i), .Q(
        \completionDataOut[1][6] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .CN(n79), .D(completionWriteData_i[5]), .E(n1255), .CP(clk_i), .Q(
        \completionDataOut[1][5] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .CN(n186), .D(completionWriteData_i[4]), .E(n1255), .CP(clk_i), .Q(
        \completionDataOut[1][4] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .CN(n41), .D(completionWriteData_i[64]), .E(n1256), .CP(clk_i), .Q(
        \completionDataOut[1][64] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .CN(n48), .D(completionWriteData_i[3]), .E(n1256), .CP(clk_i), .Q(
        \completionDataOut[1][3] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .CN(n79), .D(completionWriteData_i[2]), .E(n1256), .CP(clk_i), .Q(
        \completionDataOut[1][2] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .CN(n50), .D(completionWriteData_i[1]), .E(n1256), .CP(clk_i), .Q(
        \completionDataOut[1][1] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .CN(n77), .D(completionWriteData_i[0]), .E(n1256), .CP(clk_i), .Q(
        \completionDataOut[1][0] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .CN(n79), .D(completionWriteData_i[57]), .E(n1260), .CP(clk_i), .Q(
        \completionDataOut[1][57] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .CN(n77), .D(completionWriteData_i[56]), .E(n1258), .CP(clk_i), .Q(
        \completionDataOut[1][56] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .CN(n78), .D(completionWriteData_i[55]), .E(n1260), .CP(clk_i), .Q(
        \completionDataOut[1][55] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .CN(n186), .D(completionWriteData_i[54]), .E(n1258), .CP(clk_i), .Q(
        \completionDataOut[1][54] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .CN(n5), .D(completionWriteData_i[53]), .E(n1260), .CP(clk_i), .Q(
        \completionDataOut[1][53] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .CN(n187), .D(completionWriteData_i[52]), .E(n1258), .CP(clk_i), .Q(
        \completionDataOut[1][52] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .CN(n63), .D(completionWriteData_i[47]), .E(n1260), .CP(clk_i), .Q(
        \completionDataOut[1][47] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .CN(n80), .D(completionWriteData_i[46]), .E(n1258), .CP(clk_i), .Q(
        \completionDataOut[1][46] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .CN(n187), .D(completionWriteData_i[33]), .E(n1251), .CP(clk_i), .Q(
        \completionDataOut[1][33] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .CN(n80), .D(completionWriteData_i[32]), .E(n1251), .CP(clk_i), .Q(
        \completionDataOut[1][32] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .CN(n50), .D(completionWriteData_i[31]), .E(n1251), .CP(clk_i), .Q(
        \completionDataOut[1][31] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .CN(n63), .D(completionWriteData_i[30]), .E(n1251), .CP(clk_i), .Q(
        \completionDataOut[1][30] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .CN(n79), .D(completionWriteData_i[29]), .E(n1251), .CP(clk_i), .Q(
        \completionDataOut[1][29] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .CN(n80), .D(completionWriteData_i[28]), .E(n1251), .CP(clk_i), .Q(
        \completionDataOut[1][28] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .CN(n92), .D(completionWriteData_i[27]), .E(n1252), .CP(clk_i), .Q(
        \completionDataOut[1][27] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .CN(n48), .D(completionWriteData_i[26]), .E(n1252), .CP(clk_i), .Q(
        \completionDataOut[1][26] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .CN(n187), .D(completionWriteData_i[25]), .E(n1252), .CP(clk_i), .Q(
        \completionDataOut[1][25] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .CN(n50), .D(completionWriteData_i[24]), .E(n1252), .CP(clk_i), .Q(
        \completionDataOut[1][24] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .CN(n41), .D(completionWriteData_i[23]), .E(n1252), .CP(clk_i), .Q(
        \completionDataOut[1][23] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .CN(n41), .D(completionWriteData_i[22]), .E(n1252), .CP(clk_i), .Q(
        \completionDataOut[1][22] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .CN(n1247), .D(completionWriteData_i[66]), .E(n184), .CP(clk_i), .Q(
        \completionDataOut[0][66] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .CN(n84), .D(completionWriteData_i[65]), .E(n89), .CP(clk_i), .Q(
        \completionDataOut[0][65] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .CN(n83), .D(completionWriteData_i[56]), .E(n183), .CP(clk_i), .Q(
        \completionDataOut[0][56] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .CN(n85), .D(completionWriteData_i[54]), .E(n90), .CP(clk_i), .Q(
        \completionDataOut[0][54] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .CN(n96), .D(completionWriteData_i[47]), .E(n47), .CP(clk_i), .Q(
        \completionDataOut[0][47] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .CN(n1248), .D(completionWriteData_i[46]), .E(n89), .CP(clk_i), .Q(
        \completionDataOut[0][46] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .CN(n192), .D(completionWriteData_i[64]), .E(n90), .CP(clk_i), .Q(
        \completionDataOut[0][64] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .CN(n83), .D(completionWriteData_i[49]), .E(n182), .CP(clk_i), .Q(
        \completionDataOut[0][49] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .CN(n1247), .D(completionWriteData_i[53]), .E(n184), .CP(clk_i), .Q(
        \completionDataOut[0][53] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .CN(n85), .D(completionWriteData_i[52]), .E(n89), .CP(clk_i), .Q(
        \completionDataOut[0][52] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .CN(n191), .D(completionWriteData_i[9]), .E(n76), .CP(clk_i), .Q(
        \completionDataOut[0][9] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .CN(n193), .D(completionWriteData_i[8]), .E(n61), .CP(clk_i), .Q(
        \completionDataOut[0][8] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .CN(n71), .D(completionWriteData_i[7]), .E(n183), .CP(clk_i), .Q(
        \completionDataOut[0][7] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .CN(n86), .D(completionWriteData_i[6]), .E(n45), .CP(clk_i), .Q(
        \completionDataOut[0][6] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .CN(n1248), .D(completionWriteData_i[5]), .E(n183), .CP(clk_i), .Q(
        \completionDataOut[0][5] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .CN(n53), .D(completionWriteData_i[4]), .E(n61), .CP(clk_i), .Q(
        \completionDataOut[0][4] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .CN(n191), .D(completionWriteData_i[3]), .E(n183), .CP(clk_i), .Q(
        \completionDataOut[0][3] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .CN(n86), .D(completionWriteData_i[2]), .E(n75), .CP(clk_i), .Q(
        \completionDataOut[0][2] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .CN(n96), .D(completionWriteData_i[1]), .E(n181), .CP(clk_i), .Q(
        \completionDataOut[0][1] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .CN(n1247), .D(completionWriteData_i[0]), .E(n181), .CP(clk_i), .Q(
        \completionDataOut[0][0] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .CN(n94), .D(completionWriteData_i[33]), .E(n177), .CP(clk_i), .Q(
        \completionDataOut[4][33] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .CN(n94), .D(completionWriteData_i[32]), .E(n88), .CP(clk_i), .Q(
        \completionDataOut[4][32] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .CN(n81), .D(completionWriteData_i[27]), .E(n46), .CP(clk_i), .Q(
        \completionDataOut[4][27] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .CN(n94), .D(completionWriteData_i[26]), .E(n87), .CP(clk_i), .Q(
        \completionDataOut[4][26] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .CN(n51), .D(completionWriteData_i[22]), .E(n59), .CP(clk_i), .Q(
        \completionDataOut[4][22] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .CN(n66), .D(completionWriteData_i[21]), .E(n88), .CP(clk_i), .Q(
        \completionDataOut[4][21] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .CN(n66), .D(completionWriteData_i[20]), .E(n44), .CP(clk_i), .Q(
        \completionDataOut[4][20] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .CN(n52), .D(completionWriteData_i[16]), .E(n177), .CP(clk_i), .Q(
        \completionDataOut[4][16] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .CN(n69), .D(completionWriteData_i[14]), .E(n178), .CP(clk_i), .Q(
        \completionDataOut[4][14] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .CN(n52), .D(completionWriteData_i[10]), .E(n73), .CP(clk_i), .Q(
        \completionDataOut[4][10] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .CN(n96), .D(completionWriteData_i[63]), .E(n181), .CP(clk_i), .Q(
        \completionDataOut[0][63] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .CN(n83), .D(completionWriteData_i[62]), .E(n90), .CP(clk_i), .Q(
        \completionDataOut[0][62] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .CN(n84), .D(completionWriteData_i[61]), .E(n47), .CP(clk_i), .Q(
        \completionDataOut[0][61] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .CN(n72), .D(completionWriteData_i[60]), .E(n89), .CP(clk_i), .Q(
        \completionDataOut[0][60] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .CN(n83), .D(completionWriteData_i[59]), .E(n61), .CP(clk_i), .Q(
        \completionDataOut[0][59] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .CN(n71), .D(completionWriteData_i[58]), .E(n90), .CP(clk_i), .Q(
        \completionDataOut[0][58] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .CN(n83), .D(completionWriteData_i[39]), .E(n45), .CP(clk_i), .Q(
        \completionDataOut[0][39] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .CN(n193), .D(completionWriteData_i[38]), .E(n181), .CP(clk_i), .Q(
        \completionDataOut[0][38] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .CN(n84), .D(completionWriteData_i[37]), .E(n182), .CP(clk_i), .Q(
        \completionDataOut[0][37] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .CN(n53), .D(completionWriteData_i[36]), .E(n75), .CP(clk_i), .Q(
        \completionDataOut[0][36] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .CN(n193), .D(completionWriteData_i[35]), .E(n60), .CP(clk_i), .Q(
        \completionDataOut[0][35] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .CN(n193), .D(completionWriteData_i[34]), .E(n182), .CP(clk_i), .Q(
        \completionDataOut[0][34] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .CN(n78), .D(completionWriteData_i[63]), .E(n1262), .CP(clk_i), .Q(
        \completionDataOut[1][63] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .CN(n79), .D(completionWriteData_i[62]), .E(n1262), .CP(clk_i), .Q(
        \completionDataOut[1][62] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .CN(n41), .D(completionWriteData_i[61]), .E(n1262), .CP(clk_i), .Q(
        \completionDataOut[1][61] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .CN(n64), .D(completionWriteData_i[60]), .E(n1257), .CP(clk_i), .Q(
        \completionDataOut[1][60] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .CN(n77), .D(completionWriteData_i[59]), .E(n1259), .CP(clk_i), .Q(
        \completionDataOut[1][59] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .CN(n80), .D(completionWriteData_i[58]), .E(n1259), .CP(clk_i), .Q(
        \completionDataOut[1][58] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .CN(n190), .D(completionWriteData_i[30]), .E(n58), .CP(clk_i), .Q(
        \completionDataOut[4][30] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .CN(n190), .D(completionWriteData_i[29]), .E(n178), .CP(clk_i), .Q(
        \completionDataOut[4][29] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .CN(n42), .D(completionWriteData_i[28]), .E(n46), .CP(clk_i), .Q(
        \completionDataOut[4][28] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .CN(n67), .D(completionWriteData_i[25]), .E(n177), .CP(clk_i), .Q(
        \completionDataOut[4][25] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .CN(n93), .D(completionWriteData_i[24]), .E(n44), .CP(clk_i), .Q(
        \completionDataOut[4][24] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .CN(n93), .D(completionWriteData_i[23]), .E(n44), .CP(clk_i), .Q(
        \completionDataOut[4][23] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .CN(n67), .D(completionWriteData_i[19]), .E(n178), .CP(clk_i), .Q(
        \completionDataOut[4][19] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .CN(n3), .D(completionWriteData_i[18]), .E(n179), .CP(clk_i), .Q(
        \completionDataOut[4][18] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .CN(n82), .D(completionWriteData_i[17]), .E(n58), .CP(clk_i), .Q(
        \completionDataOut[4][17] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .CN(n69), .D(completionWriteData_i[15]), .E(n178), .CP(clk_i), .Q(
        \completionDataOut[4][15] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .CN(n93), .D(completionWriteData_i[13]), .E(n73), .CP(clk_i), .Q(
        \completionDataOut[4][13] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .CN(n190), .D(completionWriteData_i[11]), .E(n180), .CP(clk_i), .Q(
        \completionDataOut[4][11] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .CN(n42), .D(completionWriteData_i[31]), .E(n46), .CP(clk_i), .Q(
        \completionDataOut[4][31] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .CN(n82), .D(completionWriteData_i[12]), .E(n59), .CP(clk_i), .Q(
        \completionDataOut[4][12] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .CN(n66), .D(completionWriteData_i[39]), .E(n58), .CP(clk_i), .Q(
        \completionDataOut[4][39] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .CN(n81), .D(completionWriteData_i[38]), .E(n87), .CP(clk_i), .Q(
        \completionDataOut[4][38] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .CN(n67), .D(completionWriteData_i[37]), .E(n73), .CP(clk_i), .Q(
        \completionDataOut[4][37] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .CN(n81), .D(completionWriteData_i[36]), .E(n73), .CP(clk_i), .Q(
        \completionDataOut[4][36] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .CN(n81), .D(completionWriteData_i[35]), .E(n58), .CP(clk_i), .Q(
        \completionDataOut[4][35] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .CN(n52), .D(completionWriteData_i[62]), .E(n180), .CP(clk_i), .Q(
        \completionDataOut[4][62] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .CN(n51), .D(completionWriteData_i[61]), .E(n59), .CP(clk_i), .Q(
        \completionDataOut[4][61] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .CN(n94), .D(completionWriteData_i[60]), .E(n87), .CP(clk_i), .Q(
        \completionDataOut[4][60] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .CN(n42), .D(completionWriteData_i[59]), .E(n46), .CP(clk_i), .Q(
        \completionDataOut[4][59] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .CN(n68), .D(completionWriteData_i[34]), .E(n74), .CP(clk_i), .Q(
        \completionDataOut[4][34] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .CN(n51), .D(completionWriteData_i[63]), .E(n44), .CP(clk_i), .Q(
        \completionDataOut[4][63] ) );
  EDFKCNQD1 \eachCompletionReg[4].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .CN(n68), .D(completionWriteData_i[58]), .E(n74), .CP(clk_i), .Q(
        \completionDataOut[4][58] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .CN(n41), .D(completionWriteData_i[45]), .E(n1249), .CP(clk_i), .Q(
        \completionDataOut[1][45] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .CN(n187), .D(completionWriteData_i[43]), .E(n1249), .CP(clk_i), .Q(
        \completionDataOut[1][43] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .CN(n64), .D(completionWriteData_i[42]), .E(n1249), .CP(clk_i), .Q(
        \completionDataOut[1][42] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .CN(n80), .D(completionWriteData_i[41]), .E(n1249), .CP(clk_i), .Q(
        \completionDataOut[1][41] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .CN(n79), .D(completionWriteData_i[40]), .E(n1249), .CP(clk_i), .Q(
        \completionDataOut[1][40] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .CN(n48), .D(completionWriteData_i[39]), .E(n1250), .CP(clk_i), .Q(
        \completionDataOut[1][39] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .CN(n77), .D(completionWriteData_i[38]), .E(n1250), .CP(clk_i), .Q(
        \completionDataOut[1][38] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .CN(n187), .D(completionWriteData_i[37]), .E(n1250), .CP(clk_i), .Q(
        \completionDataOut[1][37] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .CN(n91), .D(completionWriteData_i[36]), .E(n1250), .CP(clk_i), .Q(
        \completionDataOut[1][36] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .CN(n64), .D(completionWriteData_i[35]), .E(n1250), .CP(clk_i), .Q(
        \completionDataOut[1][35] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .CN(n50), .D(completionWriteData_i[34]), .E(n1250), .CP(clk_i), .Q(
        \completionDataOut[1][34] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .CN(n92), .D(completionWriteData_i[21]), .E(n1253), .CP(clk_i), .Q(
        \completionDataOut[1][21] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .CN(n48), .D(completionWriteData_i[20]), .E(n1253), .CP(clk_i), .Q(
        \completionDataOut[1][20] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .CN(n186), .D(completionWriteData_i[19]), .E(n1253), .CP(clk_i), .Q(
        \completionDataOut[1][19] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .CN(n91), .D(completionWriteData_i[18]), .E(n1253), .CP(clk_i), .Q(
        \completionDataOut[1][18] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .CN(n50), .D(completionWriteData_i[17]), .E(n1253), .CP(clk_i), .Q(
        \completionDataOut[1][17] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .CN(n92), .D(completionWriteData_i[16]), .E(n1253), .CP(clk_i), .Q(
        \completionDataOut[1][16] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .CN(n91), .D(completionWriteData_i[15]), .E(n1254), .CP(clk_i), .Q(
        \completionDataOut[1][15] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .CN(n48), .D(completionWriteData_i[14]), .E(n1254), .CP(clk_i), .Q(
        \completionDataOut[1][14] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .CN(n78), .D(completionWriteData_i[13]), .E(n1254), .CP(clk_i), .Q(
        \completionDataOut[1][13] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .CN(n5), .D(completionWriteData_i[12]), .E(n1254), .CP(clk_i), .Q(
        \completionDataOut[1][12] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .CN(n63), .D(completionWriteData_i[11]), .E(n1254), .CP(clk_i), .Q(
        \completionDataOut[1][11] ) );
  EDFKCNQD1 \eachCompletionReg[1].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .CN(n78), .D(completionWriteData_i[10]), .E(n1254), .CP(clk_i), .Q(
        \completionDataOut[1][10] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .CN(n95), .D(completionWriteData_i[33]), .E(n47), .CP(clk_i), .Q(
        \completionDataOut[0][33] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .CN(n191), .D(completionWriteData_i[32]), .E(n181), .CP(clk_i), .Q(
        \completionDataOut[0][32] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .CN(n191), .D(completionWriteData_i[31]), .E(n45), .CP(clk_i), .Q(
        \completionDataOut[0][31] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .CN(n95), .D(completionWriteData_i[30]), .E(n45), .CP(clk_i), .Q(
        \completionDataOut[0][30] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .CN(n95), .D(completionWriteData_i[29]), .E(n182), .CP(clk_i), .Q(
        \completionDataOut[0][29] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .CN(n71), .D(completionWriteData_i[28]), .E(n183), .CP(clk_i), .Q(
        \completionDataOut[0][28] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .CN(n95), .D(completionWriteData_i[27]), .E(n60), .CP(clk_i), .Q(
        \completionDataOut[0][27] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .CN(n72), .D(completionWriteData_i[26]), .E(n182), .CP(clk_i), .Q(
        \completionDataOut[0][26] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .CN(n72), .D(completionWriteData_i[25]), .E(n75), .CP(clk_i), .Q(
        \completionDataOut[0][25] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .CN(n85), .D(completionWriteData_i[24]), .E(n184), .CP(clk_i), .Q(
        \completionDataOut[0][24] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .CN(n95), .D(completionWriteData_i[23]), .E(n47), .CP(clk_i), .Q(
        \completionDataOut[0][23] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .CN(n53), .D(completionWriteData_i[22]), .E(n61), .CP(clk_i), .Q(
        \completionDataOut[0][22] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .CN(n96), .D(completionWriteData_i[21]), .E(n60), .CP(clk_i), .Q(
        \completionDataOut[0][21] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .CN(n71), .D(completionWriteData_i[20]), .E(n89), .CP(clk_i), .Q(
        \completionDataOut[0][20] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .CN(n191), .D(completionWriteData_i[19]), .E(n75), .CP(clk_i), .Q(
        \completionDataOut[0][19] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .CN(n193), .D(completionWriteData_i[18]), .E(n75), .CP(clk_i), .Q(
        \completionDataOut[0][18] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .CN(n86), .D(completionWriteData_i[17]), .E(n60), .CP(clk_i), .Q(
        \completionDataOut[0][17] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .CN(n72), .D(completionWriteData_i[16]), .E(n184), .CP(clk_i), .Q(
        \completionDataOut[0][16] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .CN(n192), .D(completionWriteData_i[15]), .E(n61), .CP(clk_i), .Q(
        \completionDataOut[0][15] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .CN(n85), .D(completionWriteData_i[14]), .E(n89), .CP(clk_i), .Q(
        \completionDataOut[0][14] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .CN(n86), .D(completionWriteData_i[13]), .E(n47), .CP(clk_i), .Q(
        \completionDataOut[0][13] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .CN(n192), .D(completionWriteData_i[12]), .E(n76), .CP(clk_i), .Q(
        \completionDataOut[0][12] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .CN(n72), .D(completionWriteData_i[11]), .E(n45), .CP(clk_i), .Q(
        \completionDataOut[0][11] ) );
  EDFKCNQD1 \eachCompletionReg[0].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .CN(n86), .D(completionWriteData_i[10]), .E(n76), .CP(clk_i), .Q(
        \completionDataOut[0][10] ) );
  EDFKCNQD1 \eachManagementReg[1].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .CN(n187), .D(decodeWriteData_i[3]), .E(n176), .CP(clk_i), .Q(
        \managementDataOut[1][3] ) );
  EDFKCNQD1 \eachManagementReg[1].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .CN(n77), .D(decodeWriteData_i[2]), .E(n176), .CP(clk_i), .Q(
        \managementDataOut[1][2] ) );
  EDFKCNQD1 \eachManagementReg[1].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .CN(n92), .D(decodeWriteData_i[1]), .E(n176), .CP(clk_i), .Q(
        \managementDataOut[1][1] ) );
  EDFKCNQD1 \eachManagementReg[1].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .CN(n77), .D(decodeWriteData_i[0]), .E(n176), .CP(clk_i), .Q(
        \managementDataOut[1][0] ) );
  EDFKCNQD1 \eachManagementReg[1].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .CN(n91), .D(decodeWriteData_i[8]), .E(n509), .CP(clk_i), .Q(
        \managementDataOut[1][8] ) );
  EDFKCNQD1 \eachManagementReg[1].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .CN(n63), .D(decodeWriteData_i[7]), .E(n509), .CP(clk_i), .Q(
        \managementDataOut[1][7] ) );
  EDFKCNQD1 \eachManagementReg[1].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .CN(n91), .D(decodeWriteData_i[6]), .E(n509), .CP(clk_i), .Q(
        \managementDataOut[1][6] ) );
  EDFKCNQD1 \eachManagementReg[1].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .CN(n64), .D(decodeWriteData_i[5]), .E(n509), .CP(clk_i), .Q(
        \managementDataOut[1][5] ) );
  EDFKCNQD1 \eachManagementReg[1].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .CN(n63), .D(decodeWriteData_i[4]), .E(n509), .CP(clk_i), .Q(
        \managementDataOut[1][4] ) );
  EDFKCNQD1 \eachManagementReg[4].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .CN(n190), .D(decodeWriteData_i[7]), .E(n54), .CP(clk_i), .Q(
        \managementDataOut[4][7] ) );
  EDFKCNQD1 \eachManagementReg[4].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .CN(n189), .D(decodeWriteData_i[5]), .E(n54), .CP(clk_i), .Q(
        \managementDataOut[4][5] ) );
  EDFKCNQD1 \eachManagementReg[4].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .CN(n94), .D(decodeWriteData_i[3]), .E(n54), .CP(clk_i), .Q(
        \managementDataOut[4][3] ) );
  EDFKCNQD1 \eachManagementReg[4].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .CN(n68), .D(decodeWriteData_i[1]), .E(n321), .CP(clk_i), .Q(
        \managementDataOut[4][1] ) );
  EDFKCNQD1 \eachManagementReg[0].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .CN(n71), .D(decodeWriteData_i[4]), .E(n55), .CP(clk_i), .Q(
        \managementDataOut[0][4] ) );
  EDFKCNQD1 \eachManagementReg[0].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .CN(n193), .D(decodeWriteData_i[3]), .E(n55), .CP(clk_i), .Q(
        \managementDataOut[0][3] ) );
  EDFKCNQD1 \eachManagementReg[0].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .CN(n1248), .D(decodeWriteData_i[2]), .E(n55), .CP(clk_i), .Q(
        \managementDataOut[0][2] ) );
  EDFKCNQD1 \eachManagementReg[0].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .CN(n53), .D(decodeWriteData_i[0]), .E(n322), .CP(clk_i), .Q(
        \managementDataOut[0][0] ) );
  EDFKCNQD1 \eachManagementReg[4].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .CN(n82), .D(decodeWriteData_i[8]), .E(n321), .CP(clk_i), .Q(
        \managementDataOut[4][8] ) );
  EDFKCNQD1 \eachManagementReg[4].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .CN(n51), .D(decodeWriteData_i[6]), .E(n321), .CP(clk_i), .Q(
        \managementDataOut[4][6] ) );
  EDFKCNQD1 \eachManagementReg[0].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .CN(n72), .D(decodeWriteData_i[8]), .E(n322), .CP(clk_i), .Q(
        \managementDataOut[0][8] ) );
  EDFKCNQD1 \eachManagementReg[0].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .CN(n96), .D(decodeWriteData_i[7]), .E(n322), .CP(clk_i), .Q(
        \managementDataOut[0][7] ) );
  EDFKCNQD1 \eachManagementReg[0].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .CN(n53), .D(decodeWriteData_i[6]), .E(n322), .CP(clk_i), .Q(
        \managementDataOut[0][6] ) );
  EDFKCNQD1 \eachManagementReg[0].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .CN(n191), .D(decodeWriteData_i[5]), .E(n322), .CP(clk_i), .Q(
        \managementDataOut[0][5] ) );
  EDFKCNQD1 \eachManagementReg[0].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .CN(n71), .D(decodeWriteData_i[1]), .E(n322), .CP(clk_i), .Q(
        \managementDataOut[0][1] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[26].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][26] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[50].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][50] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[4].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[6][4] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[26].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][26] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[6].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[6][6] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[48].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][48] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[9].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[6][9] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[8].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[6][8] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[7].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[6][7] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[52].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][52] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[51].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][51] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[49].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][49] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[20].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][20] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[15].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][15] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[67].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][67] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[66].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][66] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[64].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][64] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[63].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][63] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[62].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][62] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[29].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][29] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[3].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[2][3] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[50].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][50] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[49].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][49] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[48].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][48] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[41].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][41] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[40].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][40] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[4].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[2][4] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[27].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][27] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[30].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][30] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[2].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[6][2] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[16].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][16] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[19].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][19] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[18].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][18] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[17].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][17] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[1].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[6][1] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[29].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][29] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[28].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][28] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[20].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][20] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[9].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[5][9] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[8].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[5][8] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[7].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[5][7] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[6].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[5][6] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[27].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][27] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[16].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][16] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[69].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][69] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[68].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][68] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[67].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][67] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[66].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][66] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[65].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][65] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[64].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][64] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[46].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][46] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[42].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][42] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[47].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][47] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[45].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][45] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[44].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][44] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[43].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][43] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[45].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][45] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[46].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][46] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[58].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][58] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[57].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][57] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[40].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][40] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[59].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][59] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[63].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][63] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[56].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][56] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[55].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][55] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[54].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][54] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[53].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][53] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[62].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][62] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[61].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][61] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[60].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][60] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[5].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[6][5] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[41].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][41] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[39].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][39] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[38].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][38] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[3].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[6][3] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[37].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][37] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[15].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][15] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[21].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][21] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[50].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][50] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[4].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[7][4] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[52].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][52] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[51].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][51] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[49].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][49] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[48].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][48] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[9].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[7][9] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[8].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[7][8] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[7].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[7][7] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[6].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[7][6] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[22].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][22] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[25].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][25] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[24].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][24] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[23].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][23] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[47].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][47] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[46].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][46] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[45].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][45] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[44].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][44] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[43].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][43] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[42].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][42] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[30].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][30] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[29].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][29] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[28].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][28] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[19].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][19] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[18].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][18] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[17].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][17] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[2].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[5][2] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[1].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[5][1] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[47].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][47] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[44].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][44] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[43].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][43] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[42].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][42] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[14].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][14] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[10].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][10] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[13].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][13] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[12].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][12] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[11].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][11] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[0].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[7][0] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[69].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][69] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[68].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][68] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[67].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][67] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[66].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][66] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[65].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][65] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[64].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][64] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[57].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][57] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[56].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][56] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[58].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][58] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[63].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][63] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[40].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][40] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[0].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[2][0] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[65].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][65] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[12].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][12] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[11].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][11] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[10].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][10] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[69].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][69] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[68].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][68] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[61].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][61] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[60].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][60] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[59].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][59] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[58].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][58] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[57].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][57] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[56].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][56] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[55].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][55] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[54].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][54] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[53].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][53] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[52].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][52] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[51].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][51] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[9].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[2][9] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[8].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[2][8] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[7].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[2][7] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[6].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[2][6] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[5].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[2][5] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[39].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][39] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[38].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][38] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[37].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][37] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[36].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][36] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[35].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][35] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[28].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][28] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[27].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][27] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[26].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][26] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[25].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][25] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[24].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][24] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[9].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[3][9] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[8].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[3][8] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[7].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[3][7] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[6].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[3][6] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[25].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][25] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[24].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][24] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[23].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][23] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[22].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][22] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[21].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][21] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[52].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][52] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[51].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][51] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[49].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][49] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[48].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][48] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[50].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][50] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[4].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[3][4] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[34].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][34] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[33].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][33] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[32].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][32] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[22].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][22] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[21].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][21] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[20].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][20] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[14].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][14] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[10].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][10] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[22].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][22] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[25].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][25] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[24].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][24] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[23].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][23] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[34].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][34] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[33].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][33] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[32].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][32] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[14].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][14] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[10].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][10] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[21].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][21] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[20].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][20] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[36].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][36] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[35].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][35] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[31].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][31] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[13].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][13] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[12].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][12] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[11].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[6][11] ) );
  DFQD1 \eachCompletionReg[6].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[6].completionReg/eachEnDff[0].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[6][0] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[52].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][52] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[51].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][51] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[50].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][50] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[49].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][49] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[4].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[5][4] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[48].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][48] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[55].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][55] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[54].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][54] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[53].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][53] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[62].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][62] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[61].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][61] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[60].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][60] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[5].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[5][5] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[41].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][41] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[39].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][39] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[38].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][38] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[3].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[5][3] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[59].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][59] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[37].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][37] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[14].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][14] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[13].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][13] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[11].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][11] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[10].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][10] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[0].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[3][0] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[27].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][27] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[26].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][26] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[30].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][30] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[2].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[7][2] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[16].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][16] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[19].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][19] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[18].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][18] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[17].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][17] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[15].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][15] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[1].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[7][1] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[29].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][29] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[28].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][28] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[36].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][36] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[35].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][35] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[31].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][31] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[25].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][25] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[24].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][24] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[23].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][23] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[13].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][13] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[12].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][12] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[11].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[5][11] ) );
  DFQD1 \eachCompletionReg[5].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[5].completionReg/eachEnDff[0].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[5][0] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[69].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][69] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[68].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][68] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[67].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][67] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[66].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][66] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[65].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][65] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[64].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][64] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[46].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][46] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[45].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][45] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[47].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][47] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[44].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][44] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[43].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][43] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[42].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][42] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[63].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][63] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[58].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][58] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[57].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][57] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[56].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][56] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[40].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][40] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[34].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][34] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[33].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][33] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[32].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][32] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[62].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][62] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[61].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][61] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[60].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][60] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[59].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][59] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[55].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][55] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[53].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][53] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[41].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][41] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[39].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][39] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[38].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][38] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[37].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][37] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[36].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][36] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[35].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][35] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[31].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][31] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[5].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[7][5] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[3].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[7][3] ) );
  DFQD1 \eachCompletionReg[7].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[7].completionReg/eachEnDff[54].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[7][54] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[69].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][69] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[68].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][68] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[67].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][67] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[66].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][66] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[65].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][65] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[64].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][64] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[47].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][47] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[46].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][46] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[45].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][45] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[43].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][43] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[42].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][42] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[18].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][18] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[17].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][17] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[16].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][16] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[15].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][15] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[14].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][14] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[13].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][13] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[34].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][34] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[33].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][33] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[32].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][32] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[31].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][31] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[30].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][30] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[23].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][23] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[22].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][22] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[21].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][21] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[20].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][20] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[19].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[2][19] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[2].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[2][2] ) );
  DFQD1 \eachCompletionReg[2].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[2].completionReg/eachEnDff[1].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[2][1] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[59].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][59] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[58].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][58] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[55].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][55] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[54].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][54] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[5].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[3][5] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[36].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][36] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[34].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][34] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[33].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][33] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[32].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][32] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[53].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][53] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[63].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][63] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[62].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][62] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[61].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][61] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[60].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][60] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[57].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][57] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[56].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][56] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[27].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][27] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[26].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][26] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[30].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][30] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[2].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[3][2] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[41].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][41] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[40].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][40] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[39].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][39] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[38].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][38] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[3].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[3][3] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[19].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][19] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[17].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][17] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[16].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][16] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[15].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][15] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[1].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\completionDataOut[3][1] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[29].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][29] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[28].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][28] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[18].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][18] ) );
  DFQD1 \eachManagementReg[2].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[2].managementReg/eachEnDff[3].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[2][3] ) );
  DFQD1 \eachManagementReg[2].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[2].managementReg/eachEnDff[2].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[2][2] ) );
  DFQD1 \eachManagementReg[2].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[2].managementReg/eachEnDff[1].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[2][1] ) );
  DFQD1 \eachManagementReg[2].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[2].managementReg/eachEnDff[0].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[2][0] ) );
  DFQD1 \eachManagementReg[2].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[2].managementReg/eachEnDff[8].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[2][8] ) );
  DFQD1 \eachManagementReg[2].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[2].managementReg/eachEnDff[7].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[2][7] ) );
  DFQD1 \eachManagementReg[2].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[2].managementReg/eachEnDff[6].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[2][6] ) );
  DFQD1 \eachManagementReg[2].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[2].managementReg/eachEnDff[5].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[2][5] ) );
  DFQD1 \eachManagementReg[2].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[2].managementReg/eachEnDff[4].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[2][4] ) );
  DFQD1 \eachManagementReg[5].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[5].managementReg/eachEnDff[8].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[5][8] ) );
  DFQD1 \eachManagementReg[5].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[5].managementReg/eachEnDff[0].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[5][0] ) );
  DFQD1 \eachManagementReg[5].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[5].managementReg/eachEnDff[7].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[5][7] ) );
  DFQD1 \eachManagementReg[5].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[5].managementReg/eachEnDff[1].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[5][1] ) );
  DFQD1 \eachManagementReg[7].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[7].managementReg/eachEnDff[7].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[7][7] ) );
  DFQD1 \eachManagementReg[7].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[7].managementReg/eachEnDff[3].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[7][3] ) );
  DFQD1 \eachManagementReg[7].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[7].managementReg/eachEnDff[2].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[7][2] ) );
  DFQD1 \eachManagementReg[7].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[7].managementReg/eachEnDff[0].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[7][0] ) );
  DFQD1 \eachManagementReg[6].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[6].managementReg/eachEnDff[5].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[6][5] ) );
  DFQD1 \eachManagementReg[6].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[6].managementReg/eachEnDff[4].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[6][4] ) );
  DFQD1 \eachManagementReg[6].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[6].managementReg/eachEnDff[3].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[6][3] ) );
  DFQD1 \eachManagementReg[6].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[6].managementReg/eachEnDff[2].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[6][2] ) );
  DFQD1 \eachManagementReg[7].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[7].managementReg/eachEnDff[8].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[7][8] ) );
  DFQD1 \eachManagementReg[7].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[7].managementReg/eachEnDff[6].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[7][6] ) );
  DFQD1 \eachManagementReg[7].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[7].managementReg/eachEnDff[5].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[7][5] ) );
  DFQD1 \eachManagementReg[7].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[7].managementReg/eachEnDff[4].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[7][4] ) );
  DFQD1 \eachManagementReg[7].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[7].managementReg/eachEnDff[1].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[7][1] ) );
  DFQD1 \eachManagementReg[6].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[6].managementReg/eachEnDff[8].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[6][8] ) );
  DFQD1 \eachManagementReg[6].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[6].managementReg/eachEnDff[7].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[6][7] ) );
  DFQD1 \eachManagementReg[6].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[6].managementReg/eachEnDff[6].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[6][6] ) );
  DFQD1 \eachManagementReg[6].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[6].managementReg/eachEnDff[1].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[6][1] ) );
  DFQD1 \eachManagementReg[6].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[6].managementReg/eachEnDff[0].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[6][0] ) );
  DFQD1 \eachManagementReg[3].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[3].managementReg/eachEnDff[7].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[3][7] ) );
  DFQD1 \eachManagementReg[3].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[3].managementReg/eachEnDff[3].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[3][3] ) );
  DFQD1 \eachManagementReg[3].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(\eachManagementReg[3].managementReg/eachEnDff[2].enDff/theFlop/N3 ), 
        .CP(clk_i), .Q(\managementDataOut[3][2] ) );
  EDFKCNQD2 \eachManagementReg[4].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .CN(n52), .D(decodeWriteData_i[4]), .E(n321), .CP(clk_i), .Q(
        \managementDataOut[4][4] ) );
  EDFKCNQD2 \eachManagementReg[4].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .CN(n93), .D(decodeWriteData_i[2]), .E(n321), .CP(clk_i), .Q(
        \managementDataOut[4][2] ) );
  EDFKCNQD2 \eachManagementReg[4].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .CN(n82), .D(decodeWriteData_i[0]), .E(n321), .CP(clk_i), .Q(
        \managementDataOut[4][0] ) );
  DFQD2 \eachCompletionReg[3].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[44].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][44] ) );
  EDFKCNQD4 \eachCompletionReg[1].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .CN(n48), .D(completionWriteData_i[44]), .E(n1249), .CP(clk_i), .Q(
        \completionDataOut[1][44] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[35].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][35] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[37].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][37] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[12].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][12] ) );
  DFQD1 \eachCompletionReg[3].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .D(\eachCompletionReg[3].completionReg/eachEnDff[31].enDff/theFlop/N3 ), .CP(clk_i), .Q(\completionDataOut[3][31] ) );
  CKND2D0 U1 ( .A1(n8), .A2(n9), .ZN(decodeReadData2_o[60]) );
  CKND0 U2 ( .I(n18), .ZN(n10) );
  CKND2D0 U3 ( .A1(n171), .A2(n19), .ZN(n11) );
  CKND0 U4 ( .I(n11), .ZN(n8) );
  CKND2D0 U5 ( .A1(n516), .A2(n10), .ZN(n12) );
  CKND0 U6 ( .I(n12), .ZN(n9) );
  CKND2D0 U7 ( .A1(n13), .A2(n14), .ZN(decodeReadData1_o[61]) );
  CKND0 U8 ( .I(n21), .ZN(n15) );
  CKND2D0 U9 ( .A1(n168), .A2(n22), .ZN(n16) );
  CKND0 U10 ( .I(n16), .ZN(n13) );
  CKND2D0 U11 ( .A1(n510), .A2(n15), .ZN(n17) );
  CKND0 U12 ( .I(n17), .ZN(n14) );
  IND4D2 U13 ( .A1(n20), .B1(n40), .B2(n169), .B3(n681), .ZN(
        decodeReadData1_o[44]) );
  IND4D2 U14 ( .A1(n23), .B1(n99), .B2(n531), .B3(n669), .ZN(
        decodeReadData1_o[62]) );
  CKBD1 U15 ( .I(n964), .Z(n963) );
  INVD1 U16 ( .I(n1309), .ZN(n491) );
  CKBD1 U17 ( .I(n1196), .Z(n1190) );
  CKBD1 U18 ( .I(n1196), .Z(n1188) );
  CKBD1 U19 ( .I(n1195), .Z(n1187) );
  CKBD1 U20 ( .I(n1094), .Z(n1090) );
  CKBD1 U21 ( .I(n1095), .Z(n1094) );
  CKBD1 U22 ( .I(n1093), .Z(n1092) );
  CKBD1 U23 ( .I(n1196), .Z(n1194) );
  BUFFD2 U24 ( .I(n49), .Z(n57) );
  BUFFD2 U25 ( .I(n1), .Z(n56) );
  BUFFD2 U26 ( .I(n1), .Z(n489) );
  BUFFD2 U27 ( .I(n49), .Z(n490) );
  INR2D1 U28 ( .A1(\completionDataOut[1][31] ), .B1(n116), .ZN(n114) );
  INR2D1 U29 ( .A1(\completionDataOut[3][31] ), .B1(n117), .ZN(n115) );
  INR2D1 U30 ( .A1(\completionDataOut[1][35] ), .B1(n161), .ZN(n159) );
  INR2D1 U31 ( .A1(\completionDataOut[3][35] ), .B1(n162), .ZN(n160) );
  INR2D1 U32 ( .A1(\completionDataOut[1][37] ), .B1(n161), .ZN(n157) );
  INR2D1 U33 ( .A1(\completionDataOut[3][37] ), .B1(n162), .ZN(n158) );
  AO22D0 U34 ( .A1(n1156), .A2(\completionDataOut[0][60] ), .B1(n1158), .B2(
        \completionDataOut[2][60] ), .Z(n18) );
  AOI22D1 U35 ( .A1(n1232), .A2(\completionDataOut[5][60] ), .B1(n1234), .B2(
        \completionDataOut[7][60] ), .ZN(n19) );
  AO22D0 U36 ( .A1(n1047), .A2(\completionDataOut[0][44] ), .B1(n1059), .B2(
        \completionDataOut[2][44] ), .Z(n20) );
  AO22D0 U37 ( .A1(n1055), .A2(\completionDataOut[0][61] ), .B1(n1057), .B2(
        \completionDataOut[2][61] ), .Z(n21) );
  AOI22D1 U38 ( .A1(n1130), .A2(\completionDataOut[5][61] ), .B1(n1133), .B2(
        \completionDataOut[7][61] ), .ZN(n22) );
  AO22D0 U39 ( .A1(n1055), .A2(\completionDataOut[0][62] ), .B1(n1057), .B2(
        \completionDataOut[2][62] ), .Z(n23) );
  CKBD1 U40 ( .I(n1195), .Z(n1191) );
  CKBD1 U41 ( .I(n1178), .Z(n1177) );
  CKBD1 U42 ( .I(n1093), .Z(n1091) );
  CKBD1 U43 ( .I(n1095), .Z(n1087) );
  CKBD1 U44 ( .I(n1095), .Z(n1089) );
  INVD2 U45 ( .I(decodeReadAddr1_i[2]), .ZN(n1824) );
  INVD2 U46 ( .I(n490), .ZN(n89) );
  INVD1 U47 ( .I(n62), .ZN(n187) );
  INVD1 U48 ( .I(n185), .ZN(n77) );
  INVD1 U49 ( .I(n185), .ZN(n64) );
  INVD1 U50 ( .I(n188), .ZN(n81) );
  INVD2 U51 ( .I(n489), .ZN(n87) );
  INVD2 U52 ( .I(n56), .ZN(n179) );
  INVD1 U53 ( .I(n188), .ZN(n82) );
  INVD2 U54 ( .I(n56), .ZN(n73) );
  INVD1 U55 ( .I(n65), .ZN(n94) );
  INVD2 U56 ( .I(n1), .ZN(n180) );
  INVD1 U57 ( .I(n65), .ZN(n93) );
  INVD2 U58 ( .I(n56), .ZN(n88) );
  INVD1 U59 ( .I(n188), .ZN(n67) );
  INVD2 U60 ( .I(n56), .ZN(n177) );
  INVD1 U61 ( .I(n188), .ZN(n66) );
  INVD1 U62 ( .I(n62), .ZN(n80) );
  INVD2 U63 ( .I(n57), .ZN(n183) );
  INVD1 U64 ( .I(n185), .ZN(n63) );
  INVD1 U65 ( .I(n62), .ZN(n92) );
  INVD2 U66 ( .I(n57), .ZN(n75) );
  INVD2 U67 ( .I(n49), .ZN(n184) );
  INVD2 U68 ( .I(n70), .ZN(n96) );
  INVD2 U69 ( .I(n57), .ZN(n90) );
  INVD2 U70 ( .I(n57), .ZN(n181) );
  INVD2 U71 ( .I(n490), .ZN(n60) );
  INVD2 U72 ( .I(n489), .ZN(n58) );
  INVD1 U73 ( .I(n185), .ZN(n78) );
  INVD1 U74 ( .I(n65), .ZN(n190) );
  INVD2 U75 ( .I(n489), .ZN(n59) );
  INVD2 U76 ( .I(n490), .ZN(n61) );
  INVD1 U77 ( .I(n62), .ZN(n79) );
  INVD1 U78 ( .I(n65), .ZN(n69) );
  AN2XD1 U79 ( .A1(n172), .A2(n173), .Z(n24) );
  AN2XD1 U80 ( .A1(n132), .A2(n133), .Z(n25) );
  AN2XD1 U81 ( .A1(n138), .A2(n139), .Z(n26) );
  AN2XD1 U82 ( .A1(n142), .A2(n143), .Z(n27) );
  AN2XD1 U83 ( .A1(n144), .A2(n145), .Z(n28) );
  AN2XD1 U84 ( .A1(n147), .A2(n148), .Z(n29) );
  AN2XD1 U85 ( .A1(n149), .A2(n150), .Z(n31) );
  AN2XD1 U86 ( .A1(n154), .A2(n155), .Z(n32) );
  AN2XD1 U87 ( .A1(n163), .A2(n164), .Z(n33) );
  AN2XD1 U88 ( .A1(n165), .A2(n166), .Z(n34) );
  AN2XD1 U89 ( .A1(n103), .A2(n104), .Z(n35) );
  AN2XD1 U90 ( .A1(n106), .A2(n107), .Z(n36) );
  AN2XD1 U91 ( .A1(n111), .A2(n112), .Z(n37) );
  AN2XD1 U92 ( .A1(n119), .A2(n120), .Z(n38) );
  AN2XD1 U93 ( .A1(n126), .A2(n127), .Z(n39) );
  AN2XD1 U94 ( .A1(n135), .A2(n136), .Z(n40) );
  CKBD1 U95 ( .I(n977), .Z(n966) );
  CKBD1 U96 ( .I(n1194), .Z(n1192) );
  CKBD1 U97 ( .I(n1183), .Z(n1174) );
  OR3D2 U98 ( .A1(completionWriteAddr_i[0]), .A2(n43), .A3(n1304), .Z(n1) );
  OR3D2 U99 ( .A1(completionWriteAddr_i[0]), .A2(n43), .A3(n1302), .Z(n49) );
  INVD1 U100 ( .I(n185), .ZN(n41) );
  INVD1 U101 ( .I(n188), .ZN(n42) );
  BUFFD2 U102 ( .I(resets_i[0]), .Z(n7) );
  CKBD0 U103 ( .I(completionWriteAddr_i[1]), .Z(n43) );
  INVD2 U104 ( .I(n489), .ZN(n44) );
  INVD2 U105 ( .I(n490), .ZN(n45) );
  INVD2 U106 ( .I(n56), .ZN(n46) );
  INVD2 U107 ( .I(n56), .ZN(n178) );
  INVD2 U108 ( .I(n57), .ZN(n47) );
  INVD2 U109 ( .I(n57), .ZN(n182) );
  INVD1 U110 ( .I(resets_i[1]), .ZN(n48) );
  INVD1 U111 ( .I(n62), .ZN(n186) );
  INVD1 U112 ( .I(n185), .ZN(n50) );
  INVD1 U113 ( .I(resets_i[1]), .ZN(n91) );
  INVD1 U114 ( .I(resets_i[4]), .ZN(n51) );
  INVD1 U115 ( .I(n65), .ZN(n189) );
  INVD1 U116 ( .I(resets_i[4]), .ZN(n52) );
  INVD1 U117 ( .I(n188), .ZN(n68) );
  BUFFD2 U118 ( .I(resets_i[0]), .Z(n70) );
  INVD2 U119 ( .I(n7), .ZN(n53) );
  INVD1 U120 ( .I(n70), .ZN(n192) );
  INVD1 U121 ( .I(n4), .ZN(n54) );
  OR3D2 U122 ( .A1(decodeWriteAddr_i[0]), .A2(decodeWriteAddr_i[1]), .A3(n1301), .Z(n4) );
  INVD2 U123 ( .I(n4), .ZN(n321) );
  INVD1 U124 ( .I(n174), .ZN(n55) );
  INVD2 U125 ( .I(n174), .ZN(n322) );
  INVD2 U126 ( .I(n489), .ZN(n74) );
  INVD2 U127 ( .I(n490), .ZN(n76) );
  INVD2 U128 ( .I(n5), .ZN(n62) );
  INVD2 U129 ( .I(n5), .ZN(n185) );
  INVD2 U130 ( .I(resets_i[1]), .ZN(n5) );
  INVD2 U131 ( .I(n3), .ZN(n65) );
  INVD2 U132 ( .I(n3), .ZN(n188) );
  INVD2 U133 ( .I(resets_i[4]), .ZN(n3) );
  INVD2 U134 ( .I(n7), .ZN(n71) );
  INVD2 U135 ( .I(n7), .ZN(n72) );
  INVD2 U136 ( .I(n7), .ZN(n83) );
  INVD2 U137 ( .I(n7), .ZN(n84) );
  INVD2 U138 ( .I(n7), .ZN(n193) );
  INVD2 U139 ( .I(n70), .ZN(n85) );
  INVD2 U140 ( .I(n70), .ZN(n86) );
  INVD2 U141 ( .I(n70), .ZN(n95) );
  CKBD0 U142 ( .I(n1383), .Z(n97) );
  CKBD0 U143 ( .I(n1385), .Z(n98) );
  CKBD0 U144 ( .I(n1813), .Z(n99) );
  CKBD0 U145 ( .I(n1893), .Z(n100) );
  CKBD0 U146 ( .I(n1887), .Z(n101) );
  AO22D0 U147 ( .A1(n1179), .A2(\completionDataOut[1][11] ), .B1(n1195), .B2(
        \completionDataOut[3][11] ), .Z(n1873) );
  CKND0 U148 ( .I(n1873), .ZN(n102) );
  CKND2D0 U149 ( .A1(n1178), .A2(\completionDataOut[1][8] ), .ZN(n103) );
  CKND2D0 U150 ( .A1(n1190), .A2(\completionDataOut[3][8] ), .ZN(n104) );
  CKBD0 U151 ( .I(n1846), .Z(n105) );
  CKND2D0 U152 ( .A1(n1177), .A2(\completionDataOut[1][2] ), .ZN(n106) );
  CKND2D0 U153 ( .A1(n1191), .A2(\completionDataOut[3][2] ), .ZN(n107) );
  CKBD0 U154 ( .I(n1399), .Z(n108) );
  AO22D0 U155 ( .A1(n279), .A2(\completionDataOut[1][49] ), .B1(n970), .B2(
        \completionDataOut[3][49] ), .Z(n1421) );
  CKND0 U156 ( .I(n1421), .ZN(n109) );
  CKBD0 U157 ( .I(n1423), .Z(n110) );
  CKND2D0 U158 ( .A1(n284), .A2(\completionDataOut[1][43] ), .ZN(n111) );
  CKND2D0 U159 ( .A1(n975), .A2(\completionDataOut[3][43] ), .ZN(n112) );
  BUFFD3 U160 ( .I(n979), .Z(n975) );
  CKBD0 U161 ( .I(n1463), .Z(n113) );
  NR2D1 U162 ( .A1(n114), .A2(n115), .ZN(n1481) );
  INVD1 U163 ( .I(n491), .ZN(n116) );
  CKND0 U164 ( .I(n968), .ZN(n117) );
  CKBD0 U165 ( .I(n1507), .Z(n118) );
  CKND2D0 U166 ( .A1(n282), .A2(\completionDataOut[1][19] ), .ZN(n119) );
  CKND2D0 U167 ( .A1(n977), .A2(\completionDataOut[3][19] ), .ZN(n120) );
  BUFFD3 U168 ( .I(n980), .Z(n977) );
  NR2D1 U169 ( .A1(n121), .A2(n122), .ZN(n1549) );
  INVD1 U170 ( .I(\completionDataOut[1][12] ), .ZN(n123) );
  INVD1 U171 ( .I(n963), .ZN(n124) );
  NR2D1 U172 ( .A1(n123), .A2(n124), .ZN(n121) );
  INVD1 U173 ( .I(\completionDataOut[3][12] ), .ZN(n125) );
  NR2D1 U174 ( .A1(n125), .A2(n117), .ZN(n122) );
  CKND2D0 U175 ( .A1(n285), .A2(\completionDataOut[1][7] ), .ZN(n126) );
  CKND2D0 U176 ( .A1(n978), .A2(\completionDataOut[3][7] ), .ZN(n127) );
  BUFFD3 U177 ( .I(n980), .Z(n978) );
  CKBD0 U178 ( .I(n1587), .Z(n128) );
  AO22D0 U179 ( .A1(n280), .A2(\completionDataOut[1][0] ), .B1(n965), .B2(
        \completionDataOut[3][0] ), .Z(n1589) );
  CKND0 U180 ( .I(n1589), .ZN(n129) );
  CKBD0 U181 ( .I(n1787), .Z(n130) );
  AO22D0 U182 ( .A1(n1071), .A2(\completionDataOut[1][52] ), .B1(n1093), .B2(
        \completionDataOut[3][52] ), .Z(n1781) );
  CKND0 U183 ( .I(n1781), .ZN(n131) );
  CKND2D0 U184 ( .A1(n1071), .A2(\completionDataOut[1][51] ), .ZN(n132) );
  CKND2D0 U185 ( .A1(n1092), .A2(\completionDataOut[3][51] ), .ZN(n133) );
  CKBD0 U186 ( .I(n1757), .Z(n134) );
  CKND2D0 U187 ( .A1(n1072), .A2(\completionDataOut[1][44] ), .ZN(n135) );
  CKND2D0 U188 ( .A1(n1085), .A2(\completionDataOut[3][44] ), .ZN(n136) );
  CKBD0 U189 ( .I(n1738), .Z(n137) );
  CKND2D0 U190 ( .A1(n1073), .A2(\completionDataOut[1][38] ), .ZN(n138) );
  CKND2D0 U191 ( .A1(n1091), .A2(\completionDataOut[3][38] ), .ZN(n139) );
  CKBD0 U192 ( .I(n1707), .Z(n140) );
  CKBD0 U193 ( .I(n1701), .Z(n141) );
  CKND2D0 U194 ( .A1(n1079), .A2(\completionDataOut[1][25] ), .ZN(n142) );
  CKND2D0 U195 ( .A1(n1087), .A2(\completionDataOut[3][25] ), .ZN(n143) );
  CKND2D0 U196 ( .A1(n1078), .A2(\completionDataOut[1][13] ), .ZN(n144) );
  CKND2D0 U197 ( .A1(n1094), .A2(\completionDataOut[3][13] ), .ZN(n145) );
  CKBD0 U198 ( .I(n1635), .Z(n146) );
  CKND2D0 U199 ( .A1(n1076), .A2(\completionDataOut[1][5] ), .ZN(n147) );
  CKND2D0 U200 ( .A1(n1089), .A2(\completionDataOut[3][5] ), .ZN(n148) );
  CKND2D0 U201 ( .A1(n1076), .A2(\completionDataOut[1][4] ), .ZN(n149) );
  CKND2D0 U202 ( .A1(n1090), .A2(\completionDataOut[3][4] ), .ZN(n150) );
  BUFFD3 U203 ( .I(n1077), .Z(n1076) );
  CKBD0 U204 ( .I(n2040), .Z(n151) );
  CKBD0 U205 ( .I(n2018), .Z(n152) );
  CKBD0 U206 ( .I(n2008), .Z(n153) );
  CKND2D0 U207 ( .A1(n1172), .A2(\completionDataOut[1][47] ), .ZN(n154) );
  CKND2D0 U208 ( .A1(n1194), .A2(\completionDataOut[3][47] ), .ZN(n155) );
  CKBD0 U209 ( .I(n1977), .Z(n156) );
  NR2D1 U210 ( .A1(n157), .A2(n158), .ZN(n1963) );
  NR2D1 U211 ( .A1(n159), .A2(n160), .ZN(n1957) );
  INVD1 U212 ( .I(n1174), .ZN(n161) );
  CKND0 U213 ( .I(n1192), .ZN(n162) );
  CKND2D0 U214 ( .A1(n1175), .A2(\completionDataOut[1][29] ), .ZN(n163) );
  CKND2D0 U215 ( .A1(n1187), .A2(\completionDataOut[3][29] ), .ZN(n164) );
  CKND2D0 U216 ( .A1(n1180), .A2(\completionDataOut[1][23] ), .ZN(n165) );
  CKND2D0 U217 ( .A1(n1188), .A2(\completionDataOut[3][23] ), .ZN(n166) );
  AO22D0 U218 ( .A1(n986), .A2(\completionDataOut[4][62] ), .B1(n1003), .B2(
        \completionDataOut[6][62] ), .Z(n1380) );
  CKND0 U219 ( .I(n1380), .ZN(n167) );
  CKBD0 U220 ( .I(n1812), .Z(n168) );
  CKBD0 U221 ( .I(n1755), .Z(n169) );
  CKBD0 U222 ( .I(n1666), .Z(n170) );
  CKBD0 U223 ( .I(n2041), .Z(n171) );
  CKND2D0 U224 ( .A1(n989), .A2(\completionDataOut[4][57] ), .ZN(n172) );
  CKND2D0 U225 ( .A1(n1006), .A2(\completionDataOut[6][57] ), .ZN(n173) );
  BUFFD3 U226 ( .I(n994), .Z(n989) );
  CKBD1 U227 ( .I(n30), .Z(n174) );
  INR2XD2 U228 ( .A1(n1270), .B1(resets_i[5]), .ZN(n1271) );
  CKBD0 U229 ( .I(n2060), .Z(n175) );
  OR3D0 U230 ( .A1(decodeWriteAddr_i[0]), .A2(decodeWriteAddr_i[1]), .A3(n1299), .Z(n30) );
  BUFFD2 U231 ( .I(n6), .Z(n176) );
  INVD2 U232 ( .I(n70), .ZN(n191) );
  OR2D1 U233 ( .A1(resets_i[3]), .A2(n1284), .Z(n1286) );
  AOI22D1 U234 ( .A1(n983), .A2(\completionDataOut[4][27] ), .B1(n999), .B2(
        \completionDataOut[6][27] ), .ZN(n1496) );
  AOI22D1 U235 ( .A1(n983), .A2(\completionDataOut[4][26] ), .B1(n999), .B2(
        \completionDataOut[6][26] ), .ZN(n1500) );
  AOI22D1 U236 ( .A1(n991), .A2(\completionDataOut[4][34] ), .B1(n1000), .B2(
        \completionDataOut[6][34] ), .ZN(n1470) );
  CKND1 U237 ( .I(n500), .ZN(n320) );
  AOI22D1 U238 ( .A1(n991), .A2(\completionDataOut[4][32] ), .B1(n1000), .B2(
        \completionDataOut[6][32] ), .ZN(n1478) );
  AOI22D1 U239 ( .A1(n991), .A2(\completionDataOut[4][33] ), .B1(n1000), .B2(
        \completionDataOut[6][33] ), .ZN(n1474) );
  AOI22D1 U240 ( .A1(n982), .A2(\completionDataOut[4][16] ), .B1(n998), .B2(
        \completionDataOut[6][16] ), .ZN(n1534) );
  AOI22D1 U241 ( .A1(n1018), .A2(\completionDataOut[5][64] ), .B1(n1035), .B2(
        \completionDataOut[7][64] ), .ZN(n1375) );
  AOI22D1 U242 ( .A1(n1016), .A2(\completionDataOut[5][40] ), .B1(n1033), .B2(
        \completionDataOut[7][40] ), .ZN(n1449) );
  AOI22D1 U243 ( .A1(n982), .A2(\completionDataOut[4][14] ), .B1(n998), .B2(
        \completionDataOut[6][14] ), .ZN(n1542) );
  AOI22D1 U244 ( .A1(n1015), .A2(\completionDataOut[5][27] ), .B1(n1031), .B2(
        \completionDataOut[7][27] ), .ZN(n1497) );
  AOI22D1 U245 ( .A1(n1015), .A2(\completionDataOut[5][26] ), .B1(n1031), .B2(
        \completionDataOut[7][26] ), .ZN(n1501) );
  CKBD1 U246 ( .I(n1289), .Z(n807) );
  AOI22D1 U247 ( .A1(n1023), .A2(\completionDataOut[5][34] ), .B1(n1032), .B2(
        \completionDataOut[7][34] ), .ZN(n1471) );
  AOI22D1 U248 ( .A1(n1023), .A2(\completionDataOut[5][33] ), .B1(n1032), .B2(
        \completionDataOut[7][33] ), .ZN(n1475) );
  AOI22D1 U249 ( .A1(n1023), .A2(\completionDataOut[5][32] ), .B1(n1032), .B2(
        \completionDataOut[7][32] ), .ZN(n1479) );
  AOI22D1 U250 ( .A1(n995), .A2(\completionDataOut[4][22] ), .B1(n1009), .B2(
        \completionDataOut[6][22] ), .ZN(n1514) );
  AOI22D1 U251 ( .A1(n1014), .A2(\completionDataOut[5][16] ), .B1(n1030), .B2(
        \completionDataOut[7][16] ), .ZN(n1535) );
  AOI22D1 U252 ( .A1(n995), .A2(\completionDataOut[4][20] ), .B1(n1009), .B2(
        \completionDataOut[6][20] ), .ZN(n1522) );
  INVD0 U253 ( .I(n1293), .ZN(n500) );
  AOI22D1 U254 ( .A1(n995), .A2(\completionDataOut[4][21] ), .B1(n1009), .B2(
        \completionDataOut[6][21] ), .ZN(n1518) );
  INVD1 U255 ( .I(n1294), .ZN(n507) );
  AOI22D1 U256 ( .A1(n986), .A2(\completionDataOut[4][64] ), .B1(n1003), .B2(
        \completionDataOut[6][64] ), .ZN(n1374) );
  AOI22D1 U257 ( .A1(n1022), .A2(\completionDataOut[5][46] ), .B1(n1039), .B2(
        \completionDataOut[7][46] ), .ZN(n1430) );
  AOI22D1 U258 ( .A1(n1024), .A2(\completionDataOut[5][10] ), .B1(n1042), .B2(
        \completionDataOut[7][10] ), .ZN(n1557) );
  AOI22D1 U259 ( .A1(n992), .A2(\completionDataOut[4][10] ), .B1(n1010), .B2(
        \completionDataOut[6][10] ), .ZN(n1556) );
  AOI22D1 U260 ( .A1(n1022), .A2(\completionDataOut[5][45] ), .B1(n1039), .B2(
        \completionDataOut[7][45] ), .ZN(n1434) );
  AOI22D1 U261 ( .A1(n984), .A2(\completionDataOut[4][40] ), .B1(n1001), .B2(
        \completionDataOut[6][40] ), .ZN(n1448) );
  AOI22D1 U262 ( .A1(n1014), .A2(\completionDataOut[5][14] ), .B1(n1030), .B2(
        \completionDataOut[7][14] ), .ZN(n1543) );
  AOI22D1 U263 ( .A1(n1027), .A2(\completionDataOut[5][21] ), .B1(n1041), .B2(
        \completionDataOut[7][21] ), .ZN(n1519) );
  AOI22D1 U264 ( .A1(n993), .A2(\completionDataOut[4][6] ), .B1(n1012), .B2(
        \completionDataOut[6][6] ), .ZN(n1569) );
  AOI22D1 U265 ( .A1(n1021), .A2(\completionDataOut[5][58] ), .B1(n1038), .B2(
        \completionDataOut[7][58] ), .ZN(n1393) );
  AOI22D1 U266 ( .A1(n990), .A2(\completionDataOut[4][46] ), .B1(n1007), .B2(
        \completionDataOut[6][46] ), .ZN(n1429) );
  AOI22D1 U267 ( .A1(n1027), .A2(\completionDataOut[5][22] ), .B1(n1041), .B2(
        \completionDataOut[7][22] ), .ZN(n1515) );
  INVD1 U268 ( .I(n963), .ZN(n298) );
  INVD1 U269 ( .I(n963), .ZN(n299) );
  AOI22D1 U270 ( .A1(n1027), .A2(\completionDataOut[5][20] ), .B1(n1041), .B2(
        \completionDataOut[7][20] ), .ZN(n1523) );
  INR2D1 U271 ( .A1(n1281), .B1(resets_i[2]), .ZN(n1282) );
  AOI22D1 U272 ( .A1(n1227), .A2(\completionDataOut[5][22] ), .B1(n1239), .B2(
        \completionDataOut[7][22] ), .ZN(n1913) );
  AOI22D1 U273 ( .A1(n1202), .A2(\completionDataOut[4][22] ), .B1(n1214), .B2(
        \completionDataOut[6][22] ), .ZN(n1912) );
  AOI22D1 U274 ( .A1(n1202), .A2(\completionDataOut[4][20] ), .B1(n1214), .B2(
        \completionDataOut[6][20] ), .ZN(n1904) );
  AOI22D1 U275 ( .A1(n1227), .A2(\completionDataOut[5][20] ), .B1(n1239), .B2(
        \completionDataOut[7][20] ), .ZN(n1905) );
  AOI22D1 U276 ( .A1(n1227), .A2(\completionDataOut[5][21] ), .B1(n1239), .B2(
        \completionDataOut[7][21] ), .ZN(n1909) );
  AOI22D1 U277 ( .A1(n1202), .A2(\completionDataOut[4][21] ), .B1(n1214), .B2(
        \completionDataOut[6][21] ), .ZN(n1908) );
  AOI22D1 U278 ( .A1(n1226), .A2(\completionDataOut[5][32] ), .B1(n1237), .B2(
        \completionDataOut[7][32] ), .ZN(n1947) );
  AOI22D1 U279 ( .A1(n1201), .A2(\completionDataOut[4][32] ), .B1(n1212), .B2(
        \completionDataOut[6][32] ), .ZN(n1946) );
  AOI22D1 U280 ( .A1(n1201), .A2(\completionDataOut[4][33] ), .B1(n1212), .B2(
        \completionDataOut[6][33] ), .ZN(n1950) );
  AOI22D1 U281 ( .A1(n1226), .A2(\completionDataOut[5][33] ), .B1(n1237), .B2(
        \completionDataOut[7][33] ), .ZN(n1951) );
  AOI22D1 U282 ( .A1(n1124), .A2(\completionDataOut[5][34] ), .B1(n1136), .B2(
        \completionDataOut[7][34] ), .ZN(n1723) );
  AOI22D1 U283 ( .A1(n1100), .A2(\completionDataOut[4][34] ), .B1(n1111), .B2(
        \completionDataOut[6][34] ), .ZN(n1722) );
  AOI22D1 U284 ( .A1(n1201), .A2(\completionDataOut[4][34] ), .B1(n1212), .B2(
        \completionDataOut[6][34] ), .ZN(n1954) );
  AOI22D1 U285 ( .A1(n1226), .A2(\completionDataOut[5][34] ), .B1(n1237), .B2(
        \completionDataOut[7][34] ), .ZN(n1955) );
  AOI22D1 U286 ( .A1(n1124), .A2(\completionDataOut[5][33] ), .B1(n1136), .B2(
        \completionDataOut[7][33] ), .ZN(n1719) );
  AOI22D1 U287 ( .A1(n1100), .A2(\completionDataOut[4][33] ), .B1(n1111), .B2(
        \completionDataOut[6][33] ), .ZN(n1718) );
  AOI22D1 U288 ( .A1(n1124), .A2(\completionDataOut[5][32] ), .B1(n1136), .B2(
        \completionDataOut[7][32] ), .ZN(n1715) );
  AOI22D1 U289 ( .A1(n1100), .A2(\completionDataOut[4][32] ), .B1(n1111), .B2(
        \completionDataOut[6][32] ), .ZN(n1714) );
  AOI22D1 U290 ( .A1(n1125), .A2(\completionDataOut[5][20] ), .B1(n1138), .B2(
        \completionDataOut[7][20] ), .ZN(n1674) );
  AOI22D1 U291 ( .A1(n1101), .A2(\completionDataOut[4][20] ), .B1(n1113), .B2(
        \completionDataOut[6][20] ), .ZN(n1673) );
  AOI22D1 U292 ( .A1(n1125), .A2(\completionDataOut[5][21] ), .B1(n1138), .B2(
        \completionDataOut[7][21] ), .ZN(n1678) );
  AOI22D1 U293 ( .A1(n1101), .A2(\completionDataOut[4][22] ), .B1(n1113), .B2(
        \completionDataOut[6][22] ), .ZN(n1681) );
  AOI22D1 U294 ( .A1(n1101), .A2(\completionDataOut[4][21] ), .B1(n1113), .B2(
        \completionDataOut[6][21] ), .ZN(n1677) );
  AOI22D1 U295 ( .A1(n1125), .A2(\completionDataOut[5][22] ), .B1(n1138), .B2(
        \completionDataOut[7][22] ), .ZN(n1682) );
  AOI22D1 U296 ( .A1(n989), .A2(\completionDataOut[4][58] ), .B1(n1006), .B2(
        \completionDataOut[6][58] ), .ZN(n1392) );
  OR3D1 U297 ( .A1(resets_i[6]), .A2(n1291), .A3(n1301), .Z(n1294) );
  AOI22D1 U298 ( .A1(n1224), .A2(\completionDataOut[5][45] ), .B1(n1236), .B2(
        \completionDataOut[7][45] ), .ZN(n1993) );
  AOI22D1 U299 ( .A1(n1204), .A2(\completionDataOut[4][6] ), .B1(n1215), .B2(
        \completionDataOut[6][6] ), .ZN(n1857) );
  AOI22D1 U300 ( .A1(n1098), .A2(\completionDataOut[4][42] ), .B1(n1110), .B2(
        \completionDataOut[6][42] ), .ZN(n1749) );
  AOI22D1 U301 ( .A1(n1199), .A2(\completionDataOut[4][46] ), .B1(n1211), .B2(
        \completionDataOut[6][46] ), .ZN(n1996) );
  AOI22D1 U302 ( .A1(n1224), .A2(\completionDataOut[5][46] ), .B1(n1236), .B2(
        \completionDataOut[7][46] ), .ZN(n1997) );
  AOI22D1 U303 ( .A1(n1122), .A2(\completionDataOut[5][46] ), .B1(n1135), .B2(
        \completionDataOut[7][46] ), .ZN(n1762) );
  AOI22D1 U304 ( .A1(n1230), .A2(\completionDataOut[5][16] ), .B1(n1246), .B2(
        \completionDataOut[7][16] ), .ZN(n1891) );
  AOI22D1 U305 ( .A1(n1098), .A2(\completionDataOut[4][46] ), .B1(n1110), .B2(
        \completionDataOut[6][46] ), .ZN(n1761) );
  AOI22D1 U306 ( .A1(n1205), .A2(\completionDataOut[4][16] ), .B1(n1221), .B2(
        \completionDataOut[6][16] ), .ZN(n1890) );
  AOI22D1 U307 ( .A1(n1120), .A2(\completionDataOut[5][56] ), .B1(n1134), .B2(
        \completionDataOut[7][56] ), .ZN(n1795) );
  AOI22D1 U308 ( .A1(n1230), .A2(\completionDataOut[5][14] ), .B1(n1245), .B2(
        \completionDataOut[7][14] ), .ZN(n1885) );
  AOI22D1 U309 ( .A1(n1206), .A2(\completionDataOut[4][26] ), .B1(n1213), .B2(
        \completionDataOut[6][26] ), .ZN(n1925) );
  AOI22D1 U310 ( .A1(n1199), .A2(\completionDataOut[4][42] ), .B1(n1211), .B2(
        \completionDataOut[6][42] ), .ZN(n1980) );
  AOI22D1 U311 ( .A1(n1205), .A2(\completionDataOut[4][14] ), .B1(n1220), .B2(
        \completionDataOut[6][14] ), .ZN(n1884) );
  AOI22D1 U312 ( .A1(n1231), .A2(\completionDataOut[5][26] ), .B1(n1238), .B2(
        \completionDataOut[7][26] ), .ZN(n1926) );
  AOI22D1 U313 ( .A1(n1206), .A2(\completionDataOut[4][27] ), .B1(n1213), .B2(
        \completionDataOut[6][27] ), .ZN(n1929) );
  AOI22D1 U314 ( .A1(n1231), .A2(\completionDataOut[5][27] ), .B1(n1238), .B2(
        \completionDataOut[7][27] ), .ZN(n1930) );
  AOI22D1 U315 ( .A1(n1229), .A2(\completionDataOut[5][10] ), .B1(n1240), .B2(
        \completionDataOut[7][10] ), .ZN(n1871) );
  AOI22D1 U316 ( .A1(n1204), .A2(\completionDataOut[4][10] ), .B1(n1215), .B2(
        \completionDataOut[6][10] ), .ZN(n1870) );
  AOI22D1 U317 ( .A1(n1103), .A2(\completionDataOut[4][10] ), .B1(n1114), .B2(
        \completionDataOut[6][10] ), .ZN(n1638) );
  AOI22D1 U318 ( .A1(n495), .A2(\completionDataOut[4][64] ), .B1(n1108), .B2(
        \completionDataOut[6][64] ), .ZN(n1820) );
  AOI22D1 U319 ( .A1(n1222), .A2(\completionDataOut[5][58] ), .B1(n1235), .B2(
        \completionDataOut[7][58] ), .ZN(n2038) );
  AOI22D1 U320 ( .A1(n1127), .A2(\completionDataOut[5][10] ), .B1(n1139), .B2(
        \completionDataOut[7][10] ), .ZN(n1639) );
  AOI22D1 U321 ( .A1(n1197), .A2(\completionDataOut[4][58] ), .B1(n1210), .B2(
        \completionDataOut[6][58] ), .ZN(n2037) );
  AOI22D1 U322 ( .A1(n1222), .A2(\completionDataOut[5][57] ), .B1(n1235), .B2(
        \completionDataOut[7][57] ), .ZN(n2034) );
  AOI22D1 U323 ( .A1(n1222), .A2(\completionDataOut[5][56] ), .B1(n1235), .B2(
        \completionDataOut[7][56] ), .ZN(n2030) );
  AOI22D1 U324 ( .A1(n1129), .A2(\completionDataOut[5][27] ), .B1(n1137), .B2(
        \completionDataOut[7][27] ), .ZN(n1699) );
  AOI22D1 U325 ( .A1(n1105), .A2(\completionDataOut[4][27] ), .B1(n1112), .B2(
        \completionDataOut[6][27] ), .ZN(n1698) );
  AOI22D1 U326 ( .A1(n1104), .A2(\completionDataOut[4][14] ), .B1(n1119), .B2(
        \completionDataOut[6][14] ), .ZN(n1651) );
  AOI22D1 U327 ( .A1(n1128), .A2(\completionDataOut[5][14] ), .B1(n1144), .B2(
        \completionDataOut[7][14] ), .ZN(n1652) );
  AOI22D1 U328 ( .A1(n1129), .A2(\completionDataOut[5][26] ), .B1(n1137), .B2(
        \completionDataOut[7][26] ), .ZN(n1695) );
  AOI22D1 U329 ( .A1(n1105), .A2(\completionDataOut[4][26] ), .B1(n1112), .B2(
        \completionDataOut[6][26] ), .ZN(n1694) );
  AOI22D1 U330 ( .A1(n496), .A2(\completionDataOut[4][64] ), .B1(n1209), .B2(
        \completionDataOut[6][64] ), .ZN(n2056) );
  AOI22D1 U331 ( .A1(n495), .A2(\completionDataOut[4][63] ), .B1(n1108), .B2(
        \completionDataOut[6][63] ), .ZN(n1816) );
  AOI22D1 U332 ( .A1(n1834), .A2(\completionDataOut[5][63] ), .B1(n1234), .B2(
        \completionDataOut[7][63] ), .ZN(n2053) );
  AOI22D1 U333 ( .A1(n496), .A2(\completionDataOut[4][63] ), .B1(n1209), .B2(
        \completionDataOut[6][63] ), .ZN(n2052) );
  AOI22D1 U334 ( .A1(n1132), .A2(\completionDataOut[5][63] ), .B1(n1133), .B2(
        \completionDataOut[7][63] ), .ZN(n1817) );
  CKBD1 U335 ( .I(n1248), .Z(n1247) );
  AOI22D1 U336 ( .A1(n1103), .A2(\completionDataOut[4][6] ), .B1(n1114), .B2(
        \completionDataOut[6][6] ), .ZN(n1624) );
  AOI22D1 U337 ( .A1(n1120), .A2(\completionDataOut[5][57] ), .B1(n1134), .B2(
        \completionDataOut[7][57] ), .ZN(n1799) );
  AOI22D1 U338 ( .A1(n1096), .A2(\completionDataOut[4][58] ), .B1(n1109), .B2(
        \completionDataOut[6][58] ), .ZN(n1802) );
  AOI22D1 U339 ( .A1(n1120), .A2(\completionDataOut[5][58] ), .B1(n1134), .B2(
        \completionDataOut[7][58] ), .ZN(n1803) );
  CKBD1 U340 ( .I(n944), .Z(n301) );
  CKBD1 U341 ( .I(n944), .Z(n300) );
  AOI22D1 U342 ( .A1(n994), .A2(\completionDataOut[4][42] ), .B1(n1011), .B2(
        \completionDataOut[6][42] ), .ZN(n1441) );
  OR3D1 U343 ( .A1(resets_i[6]), .A2(n1304), .A3(n1273), .Z(n1276) );
  AOI22D1 U344 ( .A1(n1200), .A2(\completionDataOut[4][40] ), .B1(n1219), .B2(
        \completionDataOut[6][40] ), .ZN(n1974) );
  AOI22D1 U345 ( .A1(n1225), .A2(\completionDataOut[5][40] ), .B1(n1244), .B2(
        \completionDataOut[7][40] ), .ZN(n1975) );
  AOI22D1 U346 ( .A1(n1099), .A2(\completionDataOut[4][40] ), .B1(n1118), .B2(
        \completionDataOut[6][40] ), .ZN(n1741) );
  AOI22D1 U347 ( .A1(n1123), .A2(\completionDataOut[5][40] ), .B1(n1143), .B2(
        \completionDataOut[7][40] ), .ZN(n1742) );
  NR2XD0 U348 ( .A1(commitReadAddr_i[2]), .A2(n1306), .ZN(n1307) );
  CKBD1 U349 ( .I(n1602), .Z(n1132) );
  NR2XD0 U350 ( .A1(commitReadAddr_i[2]), .A2(n1310), .ZN(n1311) );
  CKBD1 U351 ( .I(n1603), .Z(n1145) );
  NR2D3 U352 ( .A1(n2060), .A2(n1828), .ZN(n1834) );
  NR2D3 U353 ( .A1(n1824), .A2(n1594), .ZN(n1601) );
  OR3D0 U354 ( .A1(decodeReadAddr1_i[0]), .A2(decodeReadAddr1_i[1]), .A3(n1824), .Z(n1600) );
  OR3D0 U355 ( .A1(decodeReadAddr2_i[0]), .A2(decodeReadAddr2_i[1]), .A3(n175), 
        .Z(n1832) );
  OR3D1 U356 ( .A1(decodeReadAddr1_i[2]), .A2(decodeReadAddr1_i[0]), .A3(
        decodeReadAddr1_i[1]), .Z(n1593) );
  OR3D1 U357 ( .A1(decodeReadAddr2_i[2]), .A2(decodeReadAddr2_i[0]), .A3(
        decodeReadAddr2_i[1]), .Z(n1825) );
  AN4D1 U358 ( .A1(n1490), .A2(n1491), .A3(n1492), .A4(n1493), .Z(n2187) );
  AN4D1 U359 ( .A1(n1486), .A2(n1487), .A3(n1488), .A4(n1489), .Z(n2186) );
  AN4D1 U360 ( .A1(n1472), .A2(n1473), .A3(n1474), .A4(n1475), .Z(n2183) );
  AN4D1 U361 ( .A1(n1498), .A2(n1499), .A3(n1500), .A4(n1501), .Z(n2189) );
  AN4D1 U362 ( .A1(n1476), .A2(n1477), .A3(n1478), .A4(n1479), .Z(n2184) );
  AN4D1 U363 ( .A1(n1468), .A2(n1469), .A3(n1470), .A4(n1471), .Z(n2182) );
  AN4D1 U364 ( .A1(n1464), .A2(n1465), .A3(n1466), .A4(n1467), .Z(n2181) );
  AN4D1 U365 ( .A1(n1482), .A2(n1483), .A3(n1484), .A4(n1485), .Z(n2185) );
  AN4D1 U366 ( .A1(n1502), .A2(n1503), .A3(n1504), .A4(n1505), .Z(n2190) );
  AN4D1 U367 ( .A1(n1494), .A2(n1495), .A3(n1496), .A4(n1497), .Z(n2188) );
  AN4D1 U368 ( .A1(n1528), .A2(n1529), .A3(n1530), .A4(n1531), .Z(n2196) );
  AN4D1 U369 ( .A1(n1544), .A2(n1545), .A3(n1546), .A4(n1547), .Z(n2200) );
  AN4D1 U370 ( .A1(n1574), .A2(n1575), .A3(n1576), .A4(n1577), .Z(n2207) );
  AN4D1 U371 ( .A1(n1570), .A2(n1571), .A3(n1572), .A4(n1573), .Z(n2206) );
  AN4D1 U372 ( .A1(n1578), .A2(n1579), .A3(n1580), .A4(n1581), .Z(n2208) );
  AN4D1 U373 ( .A1(n1540), .A2(n1541), .A3(n1542), .A4(n1543), .Z(n2199) );
  AN4D1 U374 ( .A1(n1532), .A2(n1533), .A3(n1534), .A4(n1535), .Z(n2197) );
  AN4D1 U375 ( .A1(n1582), .A2(n1583), .A3(n1584), .A4(n1585), .Z(n2209) );
  AN4D1 U376 ( .A1(n1536), .A2(n1537), .A3(n1538), .A4(n1539), .Z(n2198) );
  AN4D1 U377 ( .A1(n1400), .A2(n1401), .A3(n1402), .A4(n1403), .Z(n2167) );
  AN4D1 U378 ( .A1(n1416), .A2(n1417), .A3(n1418), .A4(n1419), .Z(n2171) );
  AOI22D1 U379 ( .A1(n945), .A2(\managementDataOut[0][2] ), .B1(n958), .B2(
        \managementDataOut[2][2] ), .ZN(n1340) );
  AN4D1 U380 ( .A1(n1562), .A2(n1563), .A3(n1564), .A4(n1565), .Z(n2204) );
  AN4D1 U381 ( .A1(n1372), .A2(n1373), .A3(n1374), .A4(n1375), .Z(n2164) );
  AN4D1 U382 ( .A1(n1408), .A2(n1409), .A3(n1410), .A4(n1411), .Z(n2169) );
  AN4D1 U383 ( .A1(n1320), .A2(n1321), .A3(n1322), .A4(n1323), .Z(n2159) );
  AN4D1 U384 ( .A1(n1328), .A2(n1329), .A3(n1330), .A4(n1331), .Z(n2161) );
  AN4D1 U385 ( .A1(n1404), .A2(n1405), .A3(n1406), .A4(n1407), .Z(n2168) );
  CKAN2D0 U386 ( .A1(n520), .A2(n521), .Z(n519) );
  AN4D1 U387 ( .A1(n1446), .A2(n1447), .A3(n1448), .A4(n1449), .Z(n2177) );
  AN4D1 U388 ( .A1(n1412), .A2(n1413), .A3(n1414), .A4(n1415), .Z(n2170) );
  AN4D1 U389 ( .A1(n1508), .A2(n1509), .A3(n1510), .A4(n1511), .Z(n2191) );
  AN4D1 U390 ( .A1(n1567), .A2(n1568), .A3(n1569), .A4(n798), .Z(n2205) );
  CKAN2D0 U391 ( .A1(n646), .A2(n647), .Z(n645) );
  AN4D1 U392 ( .A1(n1512), .A2(n1513), .A3(n1514), .A4(n1515), .Z(n2192) );
  AN4D1 U393 ( .A1(n1324), .A2(n1325), .A3(n1326), .A4(n1327), .Z(n2160) );
  AN4D1 U394 ( .A1(n1316), .A2(n1317), .A3(n1318), .A4(n1319), .Z(n2158) );
  AN4D1 U395 ( .A1(n1525), .A2(n1526), .A3(n654), .A4(n1527), .Z(n2195) );
  CKAN2D0 U396 ( .A1(n529), .A2(n530), .Z(n528) );
  AN4D1 U397 ( .A1(n1516), .A2(n1517), .A3(n1518), .A4(n1519), .Z(n2193) );
  CKAN2D0 U398 ( .A1(n526), .A2(n527), .Z(n525) );
  AN4D1 U399 ( .A1(n1336), .A2(n1337), .A3(n1338), .A4(n1339), .Z(n2162) );
  AN4D1 U400 ( .A1(n1390), .A2(n1391), .A3(n1392), .A4(n1393), .Z(n2166) );
  AN4D1 U401 ( .A1(n1442), .A2(n1443), .A3(n1444), .A4(n1445), .Z(n2176) );
  AN4D1 U402 ( .A1(n1386), .A2(n1387), .A3(n1388), .A4(n1389), .Z(n2165) );
  AN4D1 U403 ( .A1(n1520), .A2(n1521), .A3(n1522), .A4(n1523), .Z(n2194) );
  AN4D1 U404 ( .A1(n1427), .A2(n1428), .A3(n1429), .A4(n1430), .Z(n2173) );
  AN4D1 U405 ( .A1(n1554), .A2(n1555), .A3(n1556), .A4(n1557), .Z(n2202) );
  AN4D1 U406 ( .A1(n1431), .A2(n1432), .A3(n1433), .A4(n1434), .Z(n2174) );
  AN4D1 U407 ( .A1(n1424), .A2(n1425), .A3(n1426), .A4(n308), .Z(n2172) );
  AN4D1 U408 ( .A1(n1458), .A2(n1459), .A3(n1460), .A4(n1461), .Z(n2180) );
  AN4D1 U409 ( .A1(n1450), .A2(n1451), .A3(n1452), .A4(n1453), .Z(n2178) );
  AN4D1 U410 ( .A1(n1550), .A2(n1551), .A3(n1552), .A4(n1553), .Z(n2201) );
  AN4D1 U411 ( .A1(n1454), .A2(n1455), .A3(n1456), .A4(n1457), .Z(n2179) );
  AN4D1 U412 ( .A1(n1439), .A2(n1440), .A3(n1441), .A4(n777), .Z(n2175) );
  AN4D1 U413 ( .A1(n1558), .A2(n1559), .A3(n1560), .A4(n1561), .Z(n2203) );
  CKAN2D0 U414 ( .A1(n649), .A2(n650), .Z(n648) );
  AN4D1 U415 ( .A1(n1675), .A2(n1676), .A3(n1677), .A4(n1678), .Z(n2092) );
  AN4D1 U416 ( .A1(n1671), .A2(n1672), .A3(n1673), .A4(n1674), .Z(n2093) );
  BUFFD1 U417 ( .I(n494), .Z(n910) );
  BUFFD1 U418 ( .I(n494), .Z(n912) );
  BUFFD1 U419 ( .I(n494), .Z(n911) );
  AN4D1 U420 ( .A1(n1910), .A2(n1911), .A3(n1912), .A4(n1913), .Z(n2141) );
  AN4D1 U421 ( .A1(n1944), .A2(n1945), .A3(n1946), .A4(n1947), .Z(n2133) );
  AN4D1 U422 ( .A1(n1906), .A2(n1907), .A3(n1908), .A4(n1909), .Z(n2142) );
  AN4D1 U423 ( .A1(n1902), .A2(n1903), .A3(n1904), .A4(n1905), .Z(n2143) );
  AN4D1 U424 ( .A1(n1948), .A2(n1949), .A3(n1950), .A4(n1951), .Z(n2132) );
  AN4D1 U425 ( .A1(n1952), .A2(n1953), .A3(n1954), .A4(n1955), .Z(n2131) );
  AN4D1 U426 ( .A1(n1712), .A2(n1713), .A3(n1714), .A4(n1715), .Z(n2084) );
  AN4D1 U427 ( .A1(n1716), .A2(n1717), .A3(n1718), .A4(n1719), .Z(n2083) );
  AN4D1 U428 ( .A1(n1720), .A2(n1721), .A3(n1722), .A4(n1723), .Z(n2082) );
  AN4D1 U429 ( .A1(n1679), .A2(n1680), .A3(n1681), .A4(n1682), .Z(n2091) );
  CKAN2D0 U430 ( .A1(n667), .A2(n668), .Z(n666) );
  CKAN2D0 U431 ( .A1(n658), .A2(n659), .Z(n657) );
  CKAN2D0 U432 ( .A1(n787), .A2(n788), .Z(n786) );
  CKAN2D0 U433 ( .A1(n628), .A2(n629), .Z(n627) );
  CKAN2D0 U434 ( .A1(n784), .A2(n785), .Z(n783) );
  CKAN2D0 U435 ( .A1(n664), .A2(n665), .Z(n663) );
  AN4D1 U436 ( .A1(n1994), .A2(n1995), .A3(n1996), .A4(n1997), .Z(n2122) );
  AN4D1 U437 ( .A1(n1923), .A2(n1924), .A3(n1925), .A4(n1926), .Z(n2138) );
  AN4D1 U438 ( .A1(n1868), .A2(n1869), .A3(n1870), .A4(n1871), .Z(n2150) );
  AN4D1 U439 ( .A1(n1927), .A2(n1928), .A3(n1929), .A4(n1930), .Z(n2137) );
  AN4D1 U440 ( .A1(n1978), .A2(n1979), .A3(n1980), .A4(n1981), .Z(n2126) );
  AN4D1 U441 ( .A1(n1888), .A2(n1889), .A3(n1890), .A4(n1891), .Z(n2146) );
  AN4D1 U442 ( .A1(n1882), .A2(n1883), .A3(n1884), .A4(n1885), .Z(n2147) );
  AN4D1 U443 ( .A1(n1855), .A2(n1856), .A3(n1857), .A4(n1858), .Z(n2153) );
  AN4D1 U444 ( .A1(n1759), .A2(n1760), .A3(n1761), .A4(n1762), .Z(n2074) );
  AN4D1 U445 ( .A1(n1747), .A2(n1748), .A3(n1749), .A4(n1750), .Z(n2076) );
  AN4D1 U446 ( .A1(n1636), .A2(n1637), .A3(n1638), .A4(n1639), .Z(n2101) );
  AN4D1 U447 ( .A1(n1649), .A2(n1650), .A3(n1651), .A4(n1652), .Z(n2098) );
  AN4D1 U448 ( .A1(n1657), .A2(n1658), .A3(n323), .A4(n331), .Z(n2096) );
  AN4D1 U449 ( .A1(n1692), .A2(n1693), .A3(n1694), .A4(n1695), .Z(n2088) );
  AN4D1 U450 ( .A1(n1696), .A2(n1697), .A3(n1698), .A4(n1699), .Z(n2087) );
  AN4D1 U451 ( .A1(n1622), .A2(n1623), .A3(n1624), .A4(n1625), .Z(n2104) );
  CKAN2D0 U452 ( .A1(n781), .A2(n782), .Z(n780) );
  CKAN2D0 U453 ( .A1(n802), .A2(n803), .Z(n801) );
  INVD1 U454 ( .I(n124), .ZN(n283) );
  INVD1 U455 ( .I(n299), .ZN(n275) );
  INVD1 U456 ( .I(n298), .ZN(n281) );
  CKAN2D0 U457 ( .A1(n523), .A2(n524), .Z(n522) );
  CKAN2D0 U458 ( .A1(n766), .A2(n767), .Z(n765) );
  CKAN2D0 U459 ( .A1(n760), .A2(n761), .Z(n759) );
  INVD1 U460 ( .I(n298), .ZN(n279) );
  INVD1 U461 ( .I(n116), .ZN(n284) );
  CKAN2D0 U462 ( .A1(n763), .A2(n764), .Z(n762) );
  INVD1 U463 ( .I(n124), .ZN(n285) );
  CKAN2D0 U464 ( .A1(n805), .A2(n806), .Z(n804) );
  INVD1 U465 ( .I(n299), .ZN(n276) );
  INVD1 U466 ( .I(n298), .ZN(n280) );
  CKAN2D0 U467 ( .A1(n661), .A2(n662), .Z(n660) );
  INVD1 U468 ( .I(n299), .ZN(n274) );
  CKAN2D0 U469 ( .A1(n793), .A2(n794), .Z(n792) );
  INVD1 U470 ( .I(n116), .ZN(n282) );
  CKAN2D0 U471 ( .A1(n652), .A2(n653), .Z(n651) );
  INVD1 U472 ( .I(n298), .ZN(n278) );
  BUFFD1 U473 ( .I(n876), .Z(n864) );
  AN4D1 U474 ( .A1(n1840), .A2(n1841), .A3(n1842), .A4(n1843), .Z(n2156) );
  AN4D1 U475 ( .A1(n1940), .A2(n1941), .A3(n1942), .A4(n1943), .Z(n2134) );
  AN4D1 U476 ( .A1(n1616), .A2(n1617), .A3(n1618), .A4(n1619), .Z(n2105) );
  AN4D1 U477 ( .A1(n1608), .A2(n1609), .A3(n1610), .A4(n1611), .Z(n2107) );
  AN4D1 U478 ( .A1(n1800), .A2(n1801), .A3(n1802), .A4(n1803), .Z(n2065) );
  AN4D1 U479 ( .A1(n1604), .A2(n1605), .A3(n1606), .A4(n1607), .Z(n2108) );
  BUFFD1 U480 ( .I(n834), .Z(n827) );
  CKAN2D0 U481 ( .A1(n595), .A2(n596), .Z(n594) );
  CKAN2D0 U482 ( .A1(n571), .A2(n572), .Z(n570) );
  AN4D1 U483 ( .A1(n1836), .A2(n1837), .A3(n1838), .A4(n1839), .Z(n2157) );
  AN4D1 U484 ( .A1(n1936), .A2(n1937), .A3(n1938), .A4(n1939), .Z(n2135) );
  CKAN2D0 U485 ( .A1(n568), .A2(n569), .Z(n567) );
  AN4D1 U486 ( .A1(n1898), .A2(n1899), .A3(n1900), .A4(n1901), .Z(n2144) );
  BUFFD1 U487 ( .I(n903), .Z(n891) );
  AN4D1 U488 ( .A1(n1851), .A2(n1852), .A3(n1853), .A4(n1854), .Z(n2154) );
  CKAN2D0 U489 ( .A1(n553), .A2(n554), .Z(n552) );
  CKAN2D0 U490 ( .A1(n613), .A2(n614), .Z(n612) );
  AN4D1 U491 ( .A1(n1667), .A2(n1668), .A3(n1669), .A4(n1670), .Z(n2094) );
  AN4D1 U492 ( .A1(n1708), .A2(n1709), .A3(n1710), .A4(n1711), .Z(n2085) );
  AN4D1 U493 ( .A1(n1847), .A2(n1848), .A3(n1849), .A4(n1850), .Z(n2155) );
  AN4D1 U494 ( .A1(n1894), .A2(n1895), .A3(n1896), .A4(n1897), .Z(n2145) );
  CKAN2D0 U495 ( .A1(n616), .A2(n617), .Z(n615) );
  CKAN2D0 U496 ( .A1(n601), .A2(n602), .Z(n600) );
  AN4D1 U497 ( .A1(n2035), .A2(n2036), .A3(n2037), .A4(n2038), .Z(n2113) );
  AN4D1 U498 ( .A1(n1739), .A2(n1740), .A3(n1741), .A4(n1742), .Z(n2078) );
  AN4D1 U499 ( .A1(n1702), .A2(n1703), .A3(n1704), .A4(n1705), .Z(n2086) );
  AN4D1 U500 ( .A1(n1612), .A2(n1613), .A3(n1614), .A4(n1615), .Z(n2106) );
  AN4D1 U501 ( .A1(n1661), .A2(n1662), .A3(n1663), .A4(n1664), .Z(n2095) );
  AN4D1 U502 ( .A1(n1972), .A2(n1973), .A3(n1974), .A4(n1975), .Z(n2127) );
  INVD1 U503 ( .I(n1276), .ZN(n494) );
  CKAN2D0 U504 ( .A1(n796), .A2(n797), .Z(n795) );
  CKAN2D0 U505 ( .A1(n619), .A2(n620), .Z(n618) );
  CKAN2D0 U506 ( .A1(n655), .A2(n656), .Z(n654) );
  CKAN2D0 U507 ( .A1(n790), .A2(n791), .Z(n789) );
  CKAN2D0 U508 ( .A1(n622), .A2(n623), .Z(n621) );
  CKBD1 U509 ( .I(n1004), .Z(n1008) );
  CKAN2D0 U510 ( .A1(n309), .A2(n310), .Z(n308) );
  CKAN2D0 U511 ( .A1(n775), .A2(n776), .Z(n774) );
  CKAN2D0 U512 ( .A1(n634), .A2(n635), .Z(n633) );
  CKAN2D0 U513 ( .A1(n772), .A2(n773), .Z(n771) );
  CKAN2D0 U514 ( .A1(n643), .A2(n644), .Z(n642) );
  CKAN2D0 U515 ( .A1(n631), .A2(n632), .Z(n630) );
  CKAN2D0 U516 ( .A1(n769), .A2(n770), .Z(n768) );
  CKBD1 U517 ( .I(n1010), .Z(n997) );
  AO22D0 U518 ( .A1(n1018), .A2(\completionDataOut[5][63] ), .B1(n1035), .B2(
        \completionDataOut[7][63] ), .Z(n1378) );
  AO22D0 U519 ( .A1(n1018), .A2(\completionDataOut[5][62] ), .B1(n1035), .B2(
        \completionDataOut[7][62] ), .Z(n1381) );
  AN4D1 U520 ( .A1(n1344), .A2(n1345), .A3(n1346), .A4(n1347), .Z(n2163) );
  CKBD1 U521 ( .I(n1009), .Z(n998) );
  BUFFD1 U522 ( .I(n929), .Z(n917) );
  AN4D1 U523 ( .A1(n2013), .A2(n2014), .A3(n2015), .A4(n2016), .Z(n2118) );
  CKAN2D0 U524 ( .A1(n541), .A2(n542), .Z(n540) );
  AN4D1 U525 ( .A1(n1818), .A2(n1819), .A3(n1820), .A4(n330), .Z(n2061) );
  AN4D1 U526 ( .A1(n1814), .A2(n1815), .A3(n1816), .A4(n1817), .Z(n2062) );
  CKAN2D0 U527 ( .A1(n538), .A2(n539), .Z(n537) );
  AN4D1 U528 ( .A1(n1775), .A2(n1776), .A3(n1777), .A4(n1778), .Z(n2070) );
  AN4D1 U529 ( .A1(n2054), .A2(n2055), .A3(n2056), .A4(n332), .Z(n2109) );
  AN4D1 U530 ( .A1(n1792), .A2(n1793), .A3(n1794), .A4(n1795), .Z(n2067) );
  AN4D1 U531 ( .A1(n2027), .A2(n2028), .A3(n2029), .A4(n2030), .Z(n2115) );
  AN4D1 U532 ( .A1(n1796), .A2(n1797), .A3(n1798), .A4(n1799), .Z(n2066) );
  AN4D1 U533 ( .A1(n2050), .A2(n2051), .A3(n2052), .A4(n2053), .Z(n2110) );
  AN4D1 U534 ( .A1(n2031), .A2(n2032), .A3(n2033), .A4(n2034), .Z(n2114) );
  CKAN2D0 U535 ( .A1(n559), .A2(n560), .Z(n558) );
  AN4D1 U536 ( .A1(n1687), .A2(n1688), .A3(n1689), .A4(n1690), .Z(n2089) );
  AN4D1 U537 ( .A1(n1683), .A2(n1684), .A3(n1685), .A4(n1686), .Z(n2090) );
  AN4D1 U538 ( .A1(n1743), .A2(n1744), .A3(n1745), .A4(n1746), .Z(n2077) );
  CKAN2D0 U539 ( .A1(n562), .A2(n563), .Z(n561) );
  AN4D1 U540 ( .A1(n1644), .A2(n1645), .A3(n1646), .A4(n1647), .Z(n2099) );
  AN4D1 U541 ( .A1(n1751), .A2(n1752), .A3(n1753), .A4(n1754), .Z(n2075) );
  AN4D1 U542 ( .A1(n1640), .A2(n1641), .A3(n1642), .A4(n1643), .Z(n2100) );
  CKAN2D0 U543 ( .A1(n544), .A2(n545), .Z(n543) );
  CKAN2D0 U544 ( .A1(n565), .A2(n566), .Z(n564) );
  AN4D1 U545 ( .A1(n1763), .A2(n1764), .A3(n1765), .A4(n1766), .Z(n2073) );
  BUFFD1 U546 ( .I(n890), .Z(n883) );
  AN4D1 U547 ( .A1(n1630), .A2(n1631), .A3(n1632), .A4(n1633), .Z(n2102) );
  BUFFD1 U548 ( .I(n890), .Z(n884) );
  AN4D1 U549 ( .A1(n1767), .A2(n1768), .A3(n1769), .A4(n1770), .Z(n2072) );
  BUFFD1 U550 ( .I(n890), .Z(n885) );
  AN4D1 U551 ( .A1(n1626), .A2(n1627), .A3(n1628), .A4(n1629), .Z(n2103) );
  AN4D1 U552 ( .A1(n1771), .A2(n1772), .A3(n1773), .A4(n1774), .Z(n2071) );
  AN4D1 U553 ( .A1(n1864), .A2(n1865), .A3(n1866), .A4(n1867), .Z(n2151) );
  AN4D1 U554 ( .A1(n1982), .A2(n1983), .A3(n1984), .A4(n1985), .Z(n2125) );
  CKAN2D0 U555 ( .A1(n598), .A2(n599), .Z(n597) );
  AN4D1 U556 ( .A1(n1986), .A2(n1987), .A3(n1988), .A4(n1989), .Z(n2124) );
  BUFFD1 U557 ( .I(n821), .Z(n812) );
  CKAN2D0 U558 ( .A1(n586), .A2(n587), .Z(n585) );
  AN4D1 U559 ( .A1(n2003), .A2(n2004), .A3(n2005), .A4(n2006), .Z(n2120) );
  AN4D1 U560 ( .A1(n1999), .A2(n2000), .A3(n2001), .A4(n2002), .Z(n2121) );
  AN4D1 U561 ( .A1(n1990), .A2(n1991), .A3(n1992), .A4(n1993), .Z(n2123) );
  CKAN2D0 U562 ( .A1(n610), .A2(n611), .Z(n609) );
  AN4D1 U563 ( .A1(n1915), .A2(n1916), .A3(n1917), .A4(n1918), .Z(n2140) );
  CKAN2D0 U564 ( .A1(n580), .A2(n581), .Z(n579) );
  AN4D1 U565 ( .A1(n1874), .A2(n1875), .A3(n1876), .A4(n1877), .Z(n2149) );
  AN4D1 U566 ( .A1(n1878), .A2(n1879), .A3(n1880), .A4(n1881), .Z(n2148) );
  AN4D1 U567 ( .A1(n2009), .A2(n2010), .A3(n2011), .A4(n2012), .Z(n2119) );
  CKAN2D0 U568 ( .A1(n607), .A2(n608), .Z(n606) );
  CKAN2D0 U569 ( .A1(n583), .A2(n584), .Z(n582) );
  BUFFD1 U570 ( .I(n821), .Z(n811) );
  AN4D1 U571 ( .A1(n1859), .A2(n1860), .A3(n1861), .A4(n1862), .Z(n2152) );
  AN4D1 U572 ( .A1(n1919), .A2(n1920), .A3(n1921), .A4(n1922), .Z(n2139) );
  CKAN2D0 U573 ( .A1(n640), .A2(n641), .Z(n639) );
  CKAN2D0 U574 ( .A1(n637), .A2(n638), .Z(n636) );
  CKBD1 U575 ( .I(n973), .Z(n971) );
  AO22D0 U576 ( .A1(n1022), .A2(\completionDataOut[5][44] ), .B1(n1043), .B2(
        \completionDataOut[7][44] ), .Z(n1437) );
  CKBD1 U577 ( .I(n1020), .Z(n1018) );
  AO22D0 U578 ( .A1(n1028), .A2(\managementDataOut[5][4] ), .B1(n1036), .B2(
        \managementDataOut[7][4] ), .Z(n1335) );
  CKBD1 U579 ( .I(n1023), .Z(n1015) );
  AO22D0 U580 ( .A1(n1020), .A2(\managementDataOut[5][0] ), .B1(n1037), .B2(
        \managementDataOut[7][0] ), .Z(n1351) );
  AO22D0 U581 ( .A1(n1020), .A2(\completionDataOut[5][69] ), .B1(n1037), .B2(
        \completionDataOut[7][69] ), .Z(n1355) );
  OR2D1 U582 ( .A1(resets_i[7]), .A2(n1295), .Z(n1298) );
  AO22D0 U583 ( .A1(n1020), .A2(\completionDataOut[5][68] ), .B1(n1037), .B2(
        \completionDataOut[7][68] ), .Z(n1359) );
  OR2D1 U584 ( .A1(resets_i[5]), .A2(n1288), .Z(n1290) );
  CKAN2D0 U585 ( .A1(n799), .A2(n800), .Z(n798) );
  INVD1 U586 ( .I(n1282), .ZN(n497) );
  CKBD1 U587 ( .I(n1012), .Z(n1010) );
  INR2XD1 U588 ( .A1(n1288), .B1(resets_i[5]), .ZN(n1289) );
  CKAN2D0 U589 ( .A1(n625), .A2(n626), .Z(n624) );
  INVD1 U590 ( .I(n1285), .ZN(n501) );
  CKBD1 U591 ( .I(n1024), .Z(n1013) );
  CKND2 U592 ( .I(n508), .ZN(n509) );
  AN4D1 U593 ( .A1(n1808), .A2(n1809), .A3(n1810), .A4(n1811), .Z(n2063) );
  AN4D1 U594 ( .A1(n1804), .A2(n1805), .A3(n1806), .A4(n1807), .Z(n2064) );
  CKAN2D0 U595 ( .A1(n691), .A2(n692), .Z(n690) );
  CKAN2D0 U596 ( .A1(n532), .A2(n533), .Z(n531) );
  CKAN2D0 U597 ( .A1(n604), .A2(n605), .Z(n603) );
  CKAN2D0 U598 ( .A1(n556), .A2(n557), .Z(n555) );
  CKAN2D0 U599 ( .A1(n736), .A2(n737), .Z(n735) );
  CKAN2D0 U600 ( .A1(n547), .A2(n548), .Z(n546) );
  CKAN2D0 U601 ( .A1(n550), .A2(n551), .Z(n549) );
  AN4D1 U602 ( .A1(n1732), .A2(n1733), .A3(n1734), .A4(n1735), .Z(n2079) );
  AN4D1 U603 ( .A1(n1728), .A2(n1729), .A3(n1730), .A4(n1731), .Z(n2080) );
  AN4D1 U604 ( .A1(n1782), .A2(n1783), .A3(n1784), .A4(n1785), .Z(n2069) );
  CKAN2D0 U605 ( .A1(n535), .A2(n536), .Z(n534) );
  AN4D1 U606 ( .A1(n1724), .A2(n1725), .A3(n1726), .A4(n1727), .Z(n2081) );
  AN4D1 U607 ( .A1(n1788), .A2(n1789), .A3(n1790), .A4(n1791), .Z(n2068) );
  AN4D1 U608 ( .A1(n1931), .A2(n1932), .A3(n1933), .A4(n1934), .Z(n2136) );
  CKAN2D0 U609 ( .A1(n742), .A2(n743), .Z(n741) );
  CKAN2D0 U610 ( .A1(n589), .A2(n590), .Z(n588) );
  AO22D0 U611 ( .A1(n1104), .A2(\completionDataOut[4][16] ), .B1(n1601), .B2(
        \completionDataOut[6][16] ), .Z(n1659) );
  AN4D1 U612 ( .A1(n1964), .A2(n1965), .A3(n1966), .A4(n1967), .Z(n2129) );
  AN4D1 U613 ( .A1(n1653), .A2(n1654), .A3(n1655), .A4(n1656), .Z(n2097) );
  AN4D1 U614 ( .A1(n1968), .A2(n1969), .A3(n1970), .A4(n1971), .Z(n2128) );
  CKAN2D0 U615 ( .A1(n709), .A2(n710), .Z(n708) );
  CKBD1 U616 ( .I(n1103), .Z(n1102) );
  BUFFD1 U617 ( .I(n848), .Z(n836) );
  CKAN2D0 U618 ( .A1(n712), .A2(n713), .Z(n711) );
  AN4D1 U619 ( .A1(n2046), .A2(n2047), .A3(n2048), .A4(n2049), .Z(n2111) );
  AN4D1 U620 ( .A1(n2042), .A2(n2043), .A3(n2044), .A4(n2045), .Z(n2112) );
  CKAN2D0 U621 ( .A1(n574), .A2(n575), .Z(n573) );
  CKAN2D0 U622 ( .A1(n757), .A2(n758), .Z(n756) );
  CKBD1 U623 ( .I(n1204), .Z(n1203) );
  AN4D1 U624 ( .A1(n2023), .A2(n2024), .A3(n2025), .A4(n2026), .Z(n2116) );
  AN4D1 U625 ( .A1(n2019), .A2(n2020), .A3(n2021), .A4(n2022), .Z(n2117) );
  CKAN2D0 U626 ( .A1(n754), .A2(n755), .Z(n753) );
  CKAN2D0 U627 ( .A1(n577), .A2(n578), .Z(n576) );
  CKAN2D0 U628 ( .A1(n700), .A2(n701), .Z(n699) );
  CKAN2D0 U629 ( .A1(n592), .A2(n593), .Z(n591) );
  CKAN2D0 U630 ( .A1(n514), .A2(n515), .Z(n513) );
  AN4D1 U631 ( .A1(n1958), .A2(n1959), .A3(n1960), .A4(n1961), .Z(n2130) );
  CKBD1 U632 ( .I(n1006), .Z(n1012) );
  CKBD1 U633 ( .I(n979), .Z(n974) );
  CKBD1 U634 ( .I(n992), .Z(n981) );
  CKBD1 U635 ( .I(n491), .Z(n964) );
  CKBD1 U636 ( .I(n1019), .Z(n1022) );
  CKBD1 U637 ( .I(n988), .Z(n986) );
  CKBD1 U638 ( .I(n1005), .Z(n1003) );
  INR2XD0 U639 ( .A1(n1284), .B1(resets_i[3]), .ZN(n1285) );
  AO22D0 U640 ( .A1(n1021), .A2(\completionDataOut[5][57] ), .B1(n1038), .B2(
        \completionDataOut[7][57] ), .Z(n1395) );
  AO22D0 U641 ( .A1(n1021), .A2(\completionDataOut[5][56] ), .B1(n1038), .B2(
        \completionDataOut[7][56] ), .Z(n1397) );
  OR2D1 U642 ( .A1(resets_i[2]), .A2(n1281), .Z(n1283) );
  CKBD1 U643 ( .I(n1006), .Z(n1002) );
  AO31D1 U644 ( .A1(decodeWriteAddr_i[0]), .A2(n194), .A3(n1296), .B(
        resets_i[7]), .Z(n1297) );
  CKAN2D0 U645 ( .A1(n778), .A2(n779), .Z(n777) );
  CKBD1 U646 ( .I(n990), .Z(n984) );
  CKBD1 U647 ( .I(n991), .Z(n983) );
  CKBD1 U648 ( .I(n1019), .Z(n1020) );
  CKAN2D0 U649 ( .A1(n721), .A2(n722), .Z(n720) );
  CKAN2D0 U650 ( .A1(n703), .A2(n704), .Z(n702) );
  CKAN2D0 U651 ( .A1(n670), .A2(n671), .Z(n669) );
  CKAN2D0 U652 ( .A1(n748), .A2(n749), .Z(n747) );
  CKBD1 U653 ( .I(n1207), .Z(n1198) );
  CKAN2D0 U654 ( .A1(n718), .A2(n719), .Z(n717) );
  CKAN2D0 U655 ( .A1(n511), .A2(n512), .Z(n510) );
  CKBD1 U656 ( .I(n1207), .Z(n1199) );
  CKAN2D0 U657 ( .A1(n682), .A2(n683), .Z(n681) );
  CKBD1 U658 ( .I(n1106), .Z(n1098) );
  CKAN2D0 U659 ( .A1(n697), .A2(n698), .Z(n696) );
  CKAN2D0 U660 ( .A1(n751), .A2(n752), .Z(n750) );
  CKAN2D0 U661 ( .A1(n724), .A2(n725), .Z(n723) );
  CKAN2D0 U662 ( .A1(n679), .A2(n680), .Z(n678) );
  CKAN2D0 U663 ( .A1(n706), .A2(n707), .Z(n705) );
  CKBD1 U664 ( .I(n1106), .Z(n1097) );
  CKAN2D0 U665 ( .A1(n676), .A2(n677), .Z(n675) );
  CKAN2D0 U666 ( .A1(n517), .A2(n518), .Z(n516) );
  CKAN2D0 U667 ( .A1(n727), .A2(n728), .Z(n726) );
  CKAN2D0 U668 ( .A1(n673), .A2(n674), .Z(n672) );
  CKAN2D0 U669 ( .A1(n715), .A2(n716), .Z(n714) );
  CKAN2D0 U670 ( .A1(n739), .A2(n740), .Z(n738) );
  NR2XD1 U671 ( .A1(resets_i[6]), .A2(n1274), .ZN(n1275) );
  BUFFD1 U672 ( .I(n863), .Z(n858) );
  BUFFD1 U673 ( .I(n863), .Z(n857) );
  BUFFD1 U674 ( .I(n863), .Z(n856) );
  INVD1 U675 ( .I(n1279), .ZN(n488) );
  INVD1 U676 ( .I(n300), .ZN(n290) );
  INVD1 U677 ( .I(n301), .ZN(n294) );
  INVD1 U678 ( .I(n944), .ZN(n288) );
  INVD1 U679 ( .I(n944), .ZN(n286) );
  CKBD1 U680 ( .I(n993), .Z(n982) );
  CKBD1 U681 ( .I(n993), .Z(n992) );
  CKBD1 U682 ( .I(n1038), .Z(n1044) );
  NR2D0 U683 ( .A1(n1291), .A2(n1301), .ZN(n1292) );
  BUFFD1 U684 ( .I(n943), .Z(n938) );
  BUFFD1 U685 ( .I(n943), .Z(n937) );
  BUFFD1 U686 ( .I(n943), .Z(n936) );
  CKBD1 U687 ( .I(n1038), .Z(n1034) );
  INVD1 U688 ( .I(n301), .ZN(n296) );
  CKBD1 U689 ( .I(n989), .Z(n985) );
  INVD1 U690 ( .I(n944), .ZN(n289) );
  CKBD1 U691 ( .I(n1011), .Z(n1007) );
  CKBD1 U692 ( .I(n987), .Z(n990) );
  CKBD1 U693 ( .I(n1037), .Z(n1035) );
  AO22D0 U694 ( .A1(n1026), .A2(\completionDataOut[5][66] ), .B1(n1037), .B2(
        \completionDataOut[7][66] ), .Z(n1367) );
  INVD1 U695 ( .I(n944), .ZN(n287) );
  INVD1 U696 ( .I(n300), .ZN(n293) );
  INVD1 U697 ( .I(n301), .ZN(n297) );
  INVD1 U698 ( .I(n300), .ZN(n291) );
  INVD1 U699 ( .I(n301), .ZN(n295) );
  INVD1 U700 ( .I(n300), .ZN(n292) );
  CKAN2D0 U701 ( .A1(n685), .A2(n686), .Z(n684) );
  AO22D0 U702 ( .A1(n1128), .A2(\completionDataOut[5][16] ), .B1(n1145), .B2(
        \completionDataOut[7][16] ), .Z(n1660) );
  CKAN2D0 U703 ( .A1(n733), .A2(n734), .Z(n732) );
  CKAN2D0 U704 ( .A1(n694), .A2(n695), .Z(n693) );
  CKAN2D0 U705 ( .A1(n730), .A2(n731), .Z(n729) );
  CKAN2D0 U706 ( .A1(n745), .A2(n746), .Z(n744) );
  CKBD1 U707 ( .I(n1078), .Z(n1075) );
  AO22D0 U708 ( .A1(n1834), .A2(\completionDataOut[5][64] ), .B1(n1234), .B2(
        \completionDataOut[7][64] ), .Z(n2057) );
  AO22D0 U709 ( .A1(n1132), .A2(\completionDataOut[5][64] ), .B1(n1133), .B2(
        \completionDataOut[7][64] ), .Z(n1821) );
  CKAN2D0 U710 ( .A1(n688), .A2(n689), .Z(n687) );
  AO22D0 U711 ( .A1(n1122), .A2(\completionDataOut[5][45] ), .B1(n1135), .B2(
        \completionDataOut[7][45] ), .Z(n1758) );
  CKBD1 U712 ( .I(n1028), .Z(n1026) );
  CKBD1 U713 ( .I(n1043), .Z(n1039) );
  CKBD1 U714 ( .I(n493), .Z(n1156) );
  CKBD1 U715 ( .I(n1232), .Z(n1224) );
  CKBD1 U716 ( .I(n492), .Z(n1055) );
  CKBD1 U717 ( .I(n1130), .Z(n1122) );
  CKND2 U718 ( .I(n945), .ZN(n944) );
  AO31D1 U719 ( .A1(completionWriteAddr_i[1]), .A2(completionWriteAddr_i[0]), 
        .A3(n1278), .B(resets_i[7]), .Z(n1279) );
  CKND2 U720 ( .I(n1832), .ZN(n496) );
  CKND2 U721 ( .I(n1600), .ZN(n495) );
  CKBD1 U722 ( .I(n1118), .Z(n1117) );
  CKBD1 U723 ( .I(n1245), .Z(n1241) );
  CKBD1 U724 ( .I(n1220), .Z(n1216) );
  CKBD1 U725 ( .I(n1118), .Z(n1116) );
  CKBD1 U726 ( .I(n1144), .Z(n1140) );
  CKBD1 U727 ( .I(n1119), .Z(n1115) );
  CKBD1 U728 ( .I(n1219), .Z(n1217) );
  BUFFD1 U729 ( .I(decodeWriteAddr_i[1]), .Z(n194) );
  NR2XD0 U730 ( .A1(n1592), .A2(n1306), .ZN(n1313) );
  OR2D0 U731 ( .A1(commitReadAddr_i[2]), .A2(n1308), .Z(n1309) );
  CKBD1 U732 ( .I(n1069), .Z(n1067) );
  CKBD1 U733 ( .I(n1170), .Z(n1169) );
  CKND2 U734 ( .I(n1593), .ZN(n492) );
  CKBD1 U735 ( .I(n1095), .Z(n1093) );
  CKBD1 U736 ( .I(n1196), .Z(n1195) );
  CKBD1 U737 ( .I(n1246), .Z(n1245) );
  CKBD1 U738 ( .I(n1221), .Z(n1220) );
  CKBD1 U739 ( .I(n1170), .Z(n1168) );
  CKBD1 U740 ( .I(n1246), .Z(n1240) );
  CKBD1 U741 ( .I(n1069), .Z(n1068) );
  CKBD1 U742 ( .I(n1221), .Z(n1215) );
  CKND2 U743 ( .I(n1825), .ZN(n493) );
  NR2XD0 U744 ( .A1(n1592), .A2(n1310), .ZN(n1315) );
  BUFFD2 U745 ( .I(n2), .Z(n1262) );
  NR2XD0 U746 ( .A1(n1273), .A2(n1304), .ZN(n1274) );
  CKBD1 U747 ( .I(completionWriteData_i[13]), .Z(n208) );
  CKBD1 U748 ( .I(completionWriteData_i[12]), .Z(n207) );
  CKBD1 U749 ( .I(completionWriteData_i[6]), .Z(n201) );
  CKBD1 U750 ( .I(completionWriteData_i[57]), .Z(n252) );
  CKBD1 U751 ( .I(completionWriteData_i[63]), .Z(n258) );
  CKBD1 U752 ( .I(completionWriteData_i[7]), .Z(n202) );
  CKBD1 U753 ( .I(completionWriteData_i[11]), .Z(n206) );
  CKBD1 U754 ( .I(completionWriteData_i[10]), .Z(n205) );
  CKBD1 U755 ( .I(completionWriteData_i[8]), .Z(n203) );
  CKBD1 U756 ( .I(completionWriteData_i[9]), .Z(n204) );
  CKBD1 U757 ( .I(completionWriteData_i[5]), .Z(n200) );
  CKBD1 U758 ( .I(completionWriteData_i[4]), .Z(n199) );
  CKBD1 U759 ( .I(completionWriteData_i[3]), .Z(n198) );
  CKBD1 U760 ( .I(completionWriteData_i[2]), .Z(n197) );
  CKBD1 U761 ( .I(completionWriteData_i[1]), .Z(n196) );
  CKBD1 U762 ( .I(completionWriteData_i[56]), .Z(n251) );
  CKBD1 U763 ( .I(completionWriteData_i[0]), .Z(n195) );
  CKBD1 U764 ( .I(completionWriteData_i[54]), .Z(n249) );
  CKBD1 U765 ( .I(completionWriteData_i[28]), .Z(n223) );
  CKBD1 U766 ( .I(decodeWriteData_i[7]), .Z(n272) );
  CKBD1 U767 ( .I(completionWriteData_i[69]), .Z(n264) );
  CKBD1 U768 ( .I(completionWriteData_i[29]), .Z(n224) );
  CKBD1 U769 ( .I(completionWriteData_i[30]), .Z(n225) );
  CKBD1 U770 ( .I(completionWriteData_i[22]), .Z(n217) );
  CKBD1 U771 ( .I(decodeWriteData_i[8]), .Z(n273) );
  CKBD1 U772 ( .I(completionWriteData_i[31]), .Z(n226) );
  CKBD1 U773 ( .I(completionWriteData_i[55]), .Z(n250) );
  CKBD1 U774 ( .I(completionWriteData_i[32]), .Z(n227) );
  CKBD1 U775 ( .I(completionWriteData_i[33]), .Z(n228) );
  CKBD1 U776 ( .I(completionWriteData_i[21]), .Z(n216) );
  CKBD1 U777 ( .I(completionWriteData_i[20]), .Z(n215) );
  CKBD1 U778 ( .I(completionWriteData_i[34]), .Z(n229) );
  CKBD1 U779 ( .I(completionWriteData_i[35]), .Z(n230) );
  CKBD1 U780 ( .I(completionWriteData_i[36]), .Z(n231) );
  CKBD1 U781 ( .I(decodeWriteData_i[0]), .Z(n265) );
  CKBD1 U782 ( .I(completionWriteData_i[27]), .Z(n222) );
  CKBD1 U783 ( .I(completionWriteData_i[65]), .Z(n260) );
  CKBD1 U784 ( .I(completionWriteData_i[64]), .Z(n259) );
  CKBD1 U785 ( .I(completionWriteData_i[62]), .Z(n257) );
  CKBD1 U786 ( .I(completionWriteData_i[66]), .Z(n261) );
  CKBD1 U787 ( .I(completionWriteData_i[60]), .Z(n255) );
  CKBD1 U788 ( .I(completionWriteData_i[26]), .Z(n221) );
  CKBD1 U789 ( .I(completionWriteData_i[67]), .Z(n262) );
  CKBD1 U790 ( .I(completionWriteData_i[24]), .Z(n219) );
  CKBD1 U791 ( .I(completionWriteData_i[59]), .Z(n254) );
  CKBD1 U792 ( .I(decodeWriteData_i[1]), .Z(n266) );
  CKBD1 U793 ( .I(completionWriteData_i[25]), .Z(n220) );
  CKBD1 U794 ( .I(completionWriteData_i[58]), .Z(n253) );
  CKBD1 U795 ( .I(decodeWriteData_i[2]), .Z(n267) );
  CKBD1 U796 ( .I(completionWriteData_i[61]), .Z(n256) );
  CKBD1 U797 ( .I(completionWriteData_i[68]), .Z(n263) );
  CKBD1 U798 ( .I(completionWriteData_i[18]), .Z(n213) );
  CKBD1 U799 ( .I(decodeWriteData_i[3]), .Z(n268) );
  CKBD1 U800 ( .I(decodeWriteData_i[4]), .Z(n269) );
  CKBD1 U801 ( .I(decodeWriteData_i[5]), .Z(n270) );
  CKBD1 U802 ( .I(decodeWriteData_i[6]), .Z(n271) );
  CKBD1 U803 ( .I(completionWriteData_i[23]), .Z(n218) );
  CKBD1 U804 ( .I(completionWriteData_i[19]), .Z(n214) );
  CKBD1 U805 ( .I(completionWriteData_i[49]), .Z(n244) );
  CKBD1 U806 ( .I(completionWriteData_i[48]), .Z(n243) );
  CKBD1 U807 ( .I(completionWriteData_i[47]), .Z(n242) );
  CKBD1 U808 ( .I(completionWriteData_i[50]), .Z(n245) );
  CKBD1 U809 ( .I(completionWriteData_i[46]), .Z(n241) );
  CKBD1 U810 ( .I(completionWriteData_i[51]), .Z(n246) );
  CKBD1 U811 ( .I(completionWriteData_i[45]), .Z(n240) );
  CKBD1 U812 ( .I(completionWriteData_i[52]), .Z(n247) );
  CKBD1 U813 ( .I(completionWriteData_i[44]), .Z(n239) );
  CKBD1 U814 ( .I(completionWriteData_i[43]), .Z(n238) );
  CKBD1 U815 ( .I(completionWriteData_i[15]), .Z(n210) );
  CKBD1 U816 ( .I(completionWriteData_i[42]), .Z(n237) );
  CKBD1 U817 ( .I(completionWriteData_i[41]), .Z(n236) );
  CKBD1 U818 ( .I(completionWriteData_i[16]), .Z(n211) );
  CKBD1 U819 ( .I(completionWriteData_i[14]), .Z(n209) );
  CKBD1 U820 ( .I(completionWriteData_i[53]), .Z(n248) );
  CKBD1 U821 ( .I(completionWriteData_i[37]), .Z(n232) );
  CKBD1 U822 ( .I(completionWriteData_i[38]), .Z(n233) );
  CKBD1 U823 ( .I(completionWriteData_i[39]), .Z(n234) );
  CKBD1 U824 ( .I(completionWriteData_i[17]), .Z(n212) );
  CKBD1 U825 ( .I(completionWriteData_i[40]), .Z(n235) );
  INVD1 U826 ( .I(n299), .ZN(n277) );
  BUFFD2 U827 ( .I(n946), .Z(n945) );
  NR2D1 U828 ( .A1(n302), .A2(n303), .ZN(n1403) );
  INVD1 U829 ( .I(\completionDataOut[5][54] ), .ZN(n304) );
  INVD1 U830 ( .I(n1026), .ZN(n305) );
  NR2D1 U831 ( .A1(n304), .A2(n305), .ZN(n302) );
  INVD1 U832 ( .I(\completionDataOut[7][54] ), .ZN(n306) );
  CKND0 U833 ( .I(n1040), .ZN(n307) );
  NR2D1 U834 ( .A1(n306), .A2(n307), .ZN(n303) );
  CKND2D0 U835 ( .A1(n1022), .A2(\completionDataOut[5][47] ), .ZN(n309) );
  CKND2D0 U836 ( .A1(n1039), .A2(\completionDataOut[7][47] ), .ZN(n310) );
  INVD1 U837 ( .I(n1283), .ZN(n311) );
  INVD1 U838 ( .I(n1283), .ZN(n312) );
  INVD1 U839 ( .I(n1298), .ZN(n313) );
  INVD1 U840 ( .I(n1298), .ZN(n314) );
  INVD1 U841 ( .I(n1290), .ZN(n315) );
  INVD1 U842 ( .I(n1290), .ZN(n316) );
  INVD1 U843 ( .I(n1286), .ZN(n317) );
  INVD1 U844 ( .I(n1286), .ZN(n318) );
  INVD1 U845 ( .I(n500), .ZN(n319) );
  CKBD1 U846 ( .I(n1229), .Z(n1228) );
  CKBD1 U847 ( .I(n1036), .Z(n1040) );
  CKBD1 U848 ( .I(n1021), .Z(n1017) );
  CKBD1 U849 ( .I(n1041), .Z(n1030) );
  CKBD1 U850 ( .I(n1042), .Z(n1029) );
  CKBD1 U851 ( .I(n1143), .Z(n1142) );
  CKBD1 U852 ( .I(n1130), .Z(n1121) );
  CKBD1 U853 ( .I(n1143), .Z(n1141) );
  CKBD1 U854 ( .I(n1127), .Z(n1126) );
  CKBD1 U855 ( .I(n1232), .Z(n1223) );
  CKBD1 U856 ( .I(n1244), .Z(n1242) );
  CKBD1 U857 ( .I(n1022), .Z(n1016) );
  AOI22D2 U858 ( .A1(n986), .A2(\completionDataOut[4][63] ), .B1(n1003), .B2(
        \completionDataOut[6][63] ), .ZN(n1377) );
  CKND0 U859 ( .I(n1659), .ZN(n323) );
  CKND0 U860 ( .I(n1335), .ZN(n324) );
  CKND0 U861 ( .I(n1351), .ZN(n325) );
  CKND0 U862 ( .I(n1355), .ZN(n326) );
  CKND0 U863 ( .I(n1359), .ZN(n327) );
  CKBD0 U864 ( .I(n1363), .Z(n328) );
  CKND0 U865 ( .I(n1367), .ZN(n329) );
  AOI22D2 U866 ( .A1(n1018), .A2(\completionDataOut[5][65] ), .B1(n1035), .B2(
        \completionDataOut[7][65] ), .ZN(n1371) );
  CKND0 U867 ( .I(n1821), .ZN(n330) );
  CKND0 U868 ( .I(n1660), .ZN(n331) );
  CKND0 U869 ( .I(n2057), .ZN(n332) );
  CKND0 U870 ( .I(n1381), .ZN(n333) );
  CKND0 U871 ( .I(n1437), .ZN(n334) );
  CKND0 U872 ( .I(n1378), .ZN(n335) );
  CKND0 U873 ( .I(n1395), .ZN(n336) );
  CKND0 U874 ( .I(n1397), .ZN(n337) );
  CKND0 U875 ( .I(n1758), .ZN(n338) );
  BUFFD2 U876 ( .I(n1599), .Z(n1095) );
  BUFFD2 U877 ( .I(n1595), .Z(n1069) );
  BUFFD2 U878 ( .I(n1831), .Z(n1196) );
  BUFFD2 U879 ( .I(n1827), .Z(n1170) );
  CKND0 U880 ( .I(n2158), .ZN(commitReadData_o[78]) );
  CKND0 U881 ( .I(n2159), .ZN(commitReadData_o[77]) );
  CKND0 U882 ( .I(n2160), .ZN(commitReadData_o[76]) );
  CKND0 U883 ( .I(n2161), .ZN(commitReadData_o[75]) );
  CKND0 U884 ( .I(n2162), .ZN(commitReadData_o[73]) );
  CKND0 U885 ( .I(n2163), .ZN(commitReadData_o[71]) );
  CKND0 U886 ( .I(n2062), .ZN(decodeReadData1_o[63]) );
  CKND0 U887 ( .I(n2145), .ZN(decodeReadData2_o[18]) );
  CKND0 U888 ( .I(n2146), .ZN(decodeReadData2_o[16]) );
  CKND0 U889 ( .I(n2061), .ZN(decodeReadData1_o[64]) );
  CKND0 U890 ( .I(n2147), .ZN(decodeReadData2_o[14]) );
  CKND0 U891 ( .I(n2148), .ZN(decodeReadData2_o[13]) );
  CKND0 U892 ( .I(n2149), .ZN(decodeReadData2_o[12]) );
  CKND0 U893 ( .I(n2150), .ZN(decodeReadData2_o[10]) );
  CKND0 U894 ( .I(n2151), .ZN(decodeReadData2_o[9]) );
  CKND0 U895 ( .I(n2152), .ZN(decodeReadData2_o[7]) );
  CKND0 U896 ( .I(n2153), .ZN(decodeReadData2_o[6]) );
  CKND0 U897 ( .I(n2154), .ZN(decodeReadData2_o[5]) );
  CKND0 U898 ( .I(n2155), .ZN(decodeReadData2_o[4]) );
  CKND0 U899 ( .I(n2156), .ZN(decodeReadData2_o[1]) );
  CKND0 U900 ( .I(n2157), .ZN(decodeReadData2_o[0]) );
  CKND0 U901 ( .I(n2164), .ZN(commitReadData_o[64]) );
  CKND0 U902 ( .I(n2165), .ZN(commitReadData_o[59]) );
  CKND0 U903 ( .I(n2166), .ZN(commitReadData_o[58]) );
  CKND0 U904 ( .I(n2167), .ZN(commitReadData_o[54]) );
  CKND0 U905 ( .I(n2144), .ZN(decodeReadData2_o[19]) );
  CKND0 U906 ( .I(n2168), .ZN(commitReadData_o[53]) );
  CKND0 U907 ( .I(n2169), .ZN(commitReadData_o[52]) );
  CKND0 U908 ( .I(n2172), .ZN(commitReadData_o[47]) );
  CKND0 U909 ( .I(n2173), .ZN(commitReadData_o[46]) );
  CKND0 U910 ( .I(n2175), .ZN(commitReadData_o[42]) );
  CKND0 U911 ( .I(n2176), .ZN(commitReadData_o[41]) );
  CKND0 U912 ( .I(n2177), .ZN(commitReadData_o[40]) );
  CKND0 U913 ( .I(n2178), .ZN(commitReadData_o[39]) );
  CKND0 U914 ( .I(n2179), .ZN(commitReadData_o[38]) );
  CKND0 U915 ( .I(n2181), .ZN(commitReadData_o[35]) );
  CKND0 U916 ( .I(n2182), .ZN(commitReadData_o[34]) );
  CKND0 U917 ( .I(n2183), .ZN(commitReadData_o[33]) );
  CKND0 U918 ( .I(n2184), .ZN(commitReadData_o[32]) );
  CKND0 U919 ( .I(n2185), .ZN(commitReadData_o[30]) );
  CKND0 U920 ( .I(n2186), .ZN(commitReadData_o[29]) );
  CKND0 U921 ( .I(n2187), .ZN(commitReadData_o[28]) );
  CKND0 U922 ( .I(n2188), .ZN(commitReadData_o[27]) );
  CKND0 U923 ( .I(n2189), .ZN(commitReadData_o[26]) );
  CKND0 U924 ( .I(n2190), .ZN(commitReadData_o[25]) );
  CKND0 U925 ( .I(n2191), .ZN(commitReadData_o[23]) );
  CKND0 U926 ( .I(n2192), .ZN(commitReadData_o[22]) );
  CKND0 U927 ( .I(n2193), .ZN(commitReadData_o[21]) );
  CKND0 U928 ( .I(n2194), .ZN(commitReadData_o[20]) );
  CKND0 U929 ( .I(n2195), .ZN(commitReadData_o[18]) );
  CKND0 U930 ( .I(n2196), .ZN(commitReadData_o[17]) );
  CKND0 U931 ( .I(n2197), .ZN(commitReadData_o[16]) );
  CKND0 U932 ( .I(n2198), .ZN(commitReadData_o[15]) );
  CKND0 U933 ( .I(n2199), .ZN(commitReadData_o[14]) );
  CKND0 U934 ( .I(n2200), .ZN(commitReadData_o[13]) );
  CKND0 U935 ( .I(n2201), .ZN(commitReadData_o[11]) );
  CKND0 U936 ( .I(n2202), .ZN(commitReadData_o[10]) );
  CKND0 U937 ( .I(n2203), .ZN(commitReadData_o[9]) );
  CKND0 U938 ( .I(n2204), .ZN(commitReadData_o[8]) );
  CKND0 U939 ( .I(n2205), .ZN(commitReadData_o[6]) );
  CKND0 U940 ( .I(n2206), .ZN(commitReadData_o[5]) );
  CKND0 U941 ( .I(n2207), .ZN(commitReadData_o[4]) );
  CKND0 U942 ( .I(n2208), .ZN(commitReadData_o[3]) );
  CKND0 U943 ( .I(n2209), .ZN(commitReadData_o[2]) );
  CKND0 U944 ( .I(n2143), .ZN(decodeReadData2_o[20]) );
  CKND0 U945 ( .I(n2063), .ZN(decodeReadData1_o[60]) );
  CKND0 U946 ( .I(n2064), .ZN(decodeReadData1_o[59]) );
  CKND0 U947 ( .I(n2065), .ZN(decodeReadData1_o[58]) );
  CKND0 U948 ( .I(n2066), .ZN(decodeReadData1_o[57]) );
  CKND0 U949 ( .I(n2067), .ZN(decodeReadData1_o[56]) );
  CKND0 U950 ( .I(n2068), .ZN(decodeReadData1_o[55]) );
  CKND0 U951 ( .I(n2069), .ZN(decodeReadData1_o[53]) );
  CKND0 U952 ( .I(n2071), .ZN(decodeReadData1_o[49]) );
  CKND0 U953 ( .I(n2072), .ZN(decodeReadData1_o[48]) );
  CKND0 U954 ( .I(n2073), .ZN(decodeReadData1_o[47]) );
  CKND0 U955 ( .I(n2074), .ZN(decodeReadData1_o[46]) );
  CKND0 U956 ( .I(n2075), .ZN(decodeReadData1_o[43]) );
  CKND0 U957 ( .I(n2076), .ZN(decodeReadData1_o[42]) );
  CKND0 U958 ( .I(n2077), .ZN(decodeReadData1_o[41]) );
  CKND0 U959 ( .I(n2078), .ZN(decodeReadData1_o[40]) );
  CKND0 U960 ( .I(n2079), .ZN(decodeReadData1_o[37]) );
  CKND0 U961 ( .I(n2080), .ZN(decodeReadData1_o[36]) );
  CKND0 U962 ( .I(n2081), .ZN(decodeReadData1_o[35]) );
  CKND0 U963 ( .I(n2082), .ZN(decodeReadData1_o[34]) );
  CKND0 U964 ( .I(n2083), .ZN(decodeReadData1_o[33]) );
  CKND0 U965 ( .I(n2084), .ZN(decodeReadData1_o[32]) );
  CKND0 U966 ( .I(n2085), .ZN(decodeReadData1_o[31]) );
  CKND0 U967 ( .I(n2086), .ZN(decodeReadData1_o[29]) );
  CKND0 U968 ( .I(n2087), .ZN(decodeReadData1_o[27]) );
  CKND0 U969 ( .I(n2088), .ZN(decodeReadData1_o[26]) );
  CKND0 U970 ( .I(n2089), .ZN(decodeReadData1_o[24]) );
  CKND0 U971 ( .I(n2090), .ZN(decodeReadData1_o[23]) );
  CKND0 U972 ( .I(n2091), .ZN(decodeReadData1_o[22]) );
  CKND0 U973 ( .I(n2092), .ZN(decodeReadData1_o[21]) );
  CKND0 U974 ( .I(n2093), .ZN(decodeReadData1_o[20]) );
  CKND0 U975 ( .I(n2094), .ZN(decodeReadData1_o[19]) );
  CKND0 U976 ( .I(n2095), .ZN(decodeReadData1_o[17]) );
  CKND0 U977 ( .I(n2096), .ZN(decodeReadData1_o[16]) );
  CKND0 U978 ( .I(n2097), .ZN(decodeReadData1_o[15]) );
  CKND0 U979 ( .I(n2098), .ZN(decodeReadData1_o[14]) );
  CKND0 U980 ( .I(n2099), .ZN(decodeReadData1_o[12]) );
  CKND0 U981 ( .I(n2100), .ZN(decodeReadData1_o[11]) );
  CKND0 U982 ( .I(n2101), .ZN(decodeReadData1_o[10]) );
  CKND0 U983 ( .I(n2102), .ZN(decodeReadData1_o[8]) );
  CKND0 U984 ( .I(n2103), .ZN(decodeReadData1_o[7]) );
  CKND0 U985 ( .I(n2104), .ZN(decodeReadData1_o[6]) );
  CKND0 U986 ( .I(n2105), .ZN(decodeReadData1_o[3]) );
  CKND0 U987 ( .I(n2106), .ZN(decodeReadData1_o[2]) );
  CKND0 U988 ( .I(n2107), .ZN(decodeReadData1_o[1]) );
  CKND0 U989 ( .I(n2108), .ZN(decodeReadData1_o[0]) );
  CKND0 U990 ( .I(n2109), .ZN(decodeReadData2_o[64]) );
  CKND0 U991 ( .I(n2110), .ZN(decodeReadData2_o[63]) );
  CKND0 U992 ( .I(n2111), .ZN(decodeReadData2_o[62]) );
  CKND0 U993 ( .I(n2112), .ZN(decodeReadData2_o[61]) );
  CKND0 U994 ( .I(n2113), .ZN(decodeReadData2_o[58]) );
  CKND0 U995 ( .I(n2125), .ZN(decodeReadData2_o[43]) );
  CKND0 U996 ( .I(n2114), .ZN(decodeReadData2_o[57]) );
  CKND0 U997 ( .I(n2115), .ZN(decodeReadData2_o[56]) );
  CKND0 U998 ( .I(n2116), .ZN(decodeReadData2_o[55]) );
  CKND0 U999 ( .I(n2117), .ZN(decodeReadData2_o[54]) );
  CKND0 U1000 ( .I(n2118), .ZN(decodeReadData2_o[52]) );
  CKND0 U1001 ( .I(n2120), .ZN(decodeReadData2_o[49]) );
  CKND0 U1002 ( .I(n2121), .ZN(decodeReadData2_o[48]) );
  CKND0 U1003 ( .I(n2122), .ZN(decodeReadData2_o[46]) );
  CKND0 U1004 ( .I(n2124), .ZN(decodeReadData2_o[44]) );
  CKND0 U1005 ( .I(n2136), .ZN(decodeReadData2_o[28]) );
  CKND0 U1006 ( .I(n2126), .ZN(decodeReadData2_o[42]) );
  CKND0 U1007 ( .I(n2127), .ZN(decodeReadData2_o[40]) );
  CKND0 U1008 ( .I(n2128), .ZN(decodeReadData2_o[39]) );
  CKND0 U1009 ( .I(n2129), .ZN(decodeReadData2_o[38]) );
  CKND0 U1010 ( .I(n2130), .ZN(decodeReadData2_o[36]) );
  CKND0 U1011 ( .I(n2131), .ZN(decodeReadData2_o[34]) );
  CKND0 U1012 ( .I(n2132), .ZN(decodeReadData2_o[33]) );
  CKND0 U1013 ( .I(n2133), .ZN(decodeReadData2_o[32]) );
  CKND0 U1014 ( .I(n2134), .ZN(decodeReadData2_o[31]) );
  CKND0 U1015 ( .I(n2135), .ZN(decodeReadData2_o[30]) );
  CKND0 U1016 ( .I(n2140), .ZN(decodeReadData2_o[24]) );
  CKND0 U1017 ( .I(n2141), .ZN(decodeReadData2_o[22]) );
  CKND0 U1018 ( .I(n2142), .ZN(decodeReadData2_o[21]) );
  CKND0 U1019 ( .I(n2137), .ZN(decodeReadData2_o[27]) );
  CKND0 U1020 ( .I(n2138), .ZN(decodeReadData2_o[26]) );
  CKND0 U1021 ( .I(n2139), .ZN(decodeReadData2_o[25]) );
  CKND0 U1022 ( .I(n2180), .ZN(commitReadData_o[37]) );
  CKND0 U1023 ( .I(n2170), .ZN(commitReadData_o[51]) );
  CKND0 U1024 ( .I(n2171), .ZN(commitReadData_o[50]) );
  CKND0 U1025 ( .I(n2174), .ZN(commitReadData_o[45]) );
  CKND0 U1026 ( .I(n2070), .ZN(decodeReadData1_o[50]) );
  CKND0 U1027 ( .I(n2119), .ZN(decodeReadData2_o[51]) );
  CKND0 U1028 ( .I(n2123), .ZN(decodeReadData2_o[45]) );
  CKBD1 U1029 ( .I(n1145), .Z(n1139) );
  CKBD1 U1030 ( .I(n1145), .Z(n1144) );
  CKBD1 U1031 ( .I(n1145), .Z(n1137) );
  CKBD1 U1032 ( .I(n1145), .Z(n1143) );
  CKBD1 U1033 ( .I(n1601), .Z(n1114) );
  CKBD1 U1034 ( .I(n1601), .Z(n1119) );
  CKBD1 U1035 ( .I(n1601), .Z(n1112) );
  CKBD1 U1036 ( .I(n1601), .Z(n1118) );
  CKBD1 U1037 ( .I(n1082), .Z(n1080) );
  BUFFD2 U1038 ( .I(n1597), .Z(n1082) );
  CKBD1 U1039 ( .I(n1183), .Z(n1181) );
  BUFFD2 U1040 ( .I(n1829), .Z(n1183) );
  CKBD1 U1041 ( .I(n495), .Z(n1107) );
  CKBD1 U1042 ( .I(n495), .Z(n1099) );
  CKBD1 U1043 ( .I(n495), .Z(n1096) );
  CKBD1 U1044 ( .I(n495), .Z(n1106) );
  CKBD1 U1045 ( .I(n496), .Z(n1208) );
  CKBD1 U1046 ( .I(n496), .Z(n1200) );
  CKBD1 U1047 ( .I(n496), .Z(n1197) );
  CKBD1 U1048 ( .I(n496), .Z(n1207) );
  CKBD1 U1049 ( .I(n1132), .Z(n1131) );
  CKBD1 U1050 ( .I(n1132), .Z(n1123) );
  CKBD1 U1051 ( .I(n1132), .Z(n1120) );
  CKBD1 U1052 ( .I(n1132), .Z(n1130) );
  CKBD1 U1053 ( .I(n1834), .Z(n1233) );
  CKBD1 U1054 ( .I(n1834), .Z(n1225) );
  CKBD1 U1055 ( .I(n1834), .Z(n1222) );
  CKBD1 U1056 ( .I(n1834), .Z(n1232) );
  NR3D1 U1057 ( .A1(commitReadAddr_i[2]), .A2(commitReadAddr_i[0]), .A3(
        commitReadAddr_i[1]), .ZN(n1305) );
  NR3D1 U1058 ( .A1(commitReadAddr_i[0]), .A2(commitReadAddr_i[1]), .A3(n1592), 
        .ZN(n1312) );
  BUFFD2 U1059 ( .I(n1257), .Z(n1256) );
  BUFFD2 U1060 ( .I(n1257), .Z(n1255) );
  BUFFD2 U1061 ( .I(n1262), .Z(n1257) );
  INVD1 U1062 ( .I(commitReadAddr_i[2]), .ZN(n1592) );
  BUFFD2 U1063 ( .I(n1259), .Z(n1251) );
  BUFFD2 U1064 ( .I(n1259), .Z(n1252) );
  BUFFD2 U1065 ( .I(n1262), .Z(n1259) );
  BUFFD2 U1066 ( .I(n1261), .Z(n1260) );
  BUFFD2 U1067 ( .I(n1261), .Z(n1258) );
  BUFFD2 U1068 ( .I(n1262), .Z(n1261) );
  BUFFD2 U1069 ( .I(n1258), .Z(n1254) );
  BUFFD2 U1070 ( .I(n1258), .Z(n1253) );
  BUFFD2 U1071 ( .I(n1260), .Z(n1249) );
  BUFFD2 U1072 ( .I(n1260), .Z(n1250) );
  ND2D1 U1073 ( .A1(completionWriteEn_i), .A2(completionWriteAddr_i[2]), .ZN(
        n1304) );
  INVD1 U1074 ( .I(n497), .ZN(n498) );
  INVD1 U1075 ( .I(n497), .ZN(n499) );
  NR2D0 U1076 ( .A1(resets_i[6]), .A2(n1292), .ZN(n1293) );
  INVD1 U1077 ( .I(n501), .ZN(n502) );
  INVD1 U1078 ( .I(n501), .ZN(n503) );
  INVD1 U1079 ( .I(n1297), .ZN(n504) );
  INVD1 U1080 ( .I(n1297), .ZN(n505) );
  INVD1 U1081 ( .I(n1294), .ZN(n506) );
  INVD1 U1082 ( .I(n176), .ZN(n508) );
  CKND2D0 U1083 ( .A1(n1080), .A2(\completionDataOut[1][61] ), .ZN(n511) );
  CKND2D0 U1084 ( .A1(n1083), .A2(\completionDataOut[3][61] ), .ZN(n512) );
  CKND2D0 U1085 ( .A1(n1075), .A2(\completionDataOut[1][18] ), .ZN(n514) );
  CKND2D0 U1086 ( .A1(n1088), .A2(\completionDataOut[3][18] ), .ZN(n515) );
  CKND2D0 U1087 ( .A1(n1181), .A2(\completionDataOut[1][60] ), .ZN(n517) );
  CKND2D0 U1088 ( .A1(n1184), .A2(\completionDataOut[3][60] ), .ZN(n518) );
  CKND2D0 U1089 ( .A1(n281), .A2(\completionDataOut[1][63] ), .ZN(n520) );
  CKND2D0 U1090 ( .A1(n971), .A2(\completionDataOut[3][63] ), .ZN(n521) );
  ND4D8 U1091 ( .A1(n1376), .A2(n519), .A3(n1377), .A4(n335), .ZN(
        commitReadData_o[63]) );
  CKND2D0 U1092 ( .A1(n491), .A2(\completionDataOut[1][62] ), .ZN(n523) );
  CKND2D0 U1093 ( .A1(n971), .A2(\completionDataOut[3][62] ), .ZN(n524) );
  ND4D8 U1094 ( .A1(n1379), .A2(n522), .A3(n167), .A4(n333), .ZN(
        commitReadData_o[62]) );
  CKND2D0 U1095 ( .A1(n284), .A2(\completionDataOut[1][57] ), .ZN(n526) );
  CKND2D0 U1096 ( .A1(n974), .A2(\completionDataOut[3][57] ), .ZN(n527) );
  ND4D8 U1097 ( .A1(n1394), .A2(n525), .A3(n24), .A4(n336), .ZN(
        commitReadData_o[57]) );
  CKND2D0 U1098 ( .A1(n285), .A2(\completionDataOut[1][56] ), .ZN(n529) );
  CKND2D0 U1099 ( .A1(n974), .A2(\completionDataOut[3][56] ), .ZN(n530) );
  CKND2D0 U1100 ( .A1(n1106), .A2(\completionDataOut[4][62] ), .ZN(n532) );
  CKND2D0 U1101 ( .A1(n1108), .A2(\completionDataOut[6][62] ), .ZN(n533) );
  CKND2D0 U1102 ( .A1(n1096), .A2(\completionDataOut[4][54] ), .ZN(n535) );
  CKND2D0 U1103 ( .A1(n1109), .A2(\completionDataOut[6][54] ), .ZN(n536) );
  CKND2D0 U1104 ( .A1(n1097), .A2(\completionDataOut[4][52] ), .ZN(n538) );
  CKND2D0 U1105 ( .A1(n1118), .A2(\completionDataOut[6][52] ), .ZN(n539) );
  CKND2D0 U1106 ( .A1(n1097), .A2(\completionDataOut[4][51] ), .ZN(n541) );
  CKND2D0 U1107 ( .A1(n1117), .A2(\completionDataOut[6][51] ), .ZN(n542) );
  CKND2D0 U1108 ( .A1(n1098), .A2(\completionDataOut[4][45] ), .ZN(n544) );
  CKND2D0 U1109 ( .A1(n1110), .A2(\completionDataOut[6][45] ), .ZN(n545) );
  ND4D8 U1110 ( .A1(n1756), .A2(n134), .A3(n543), .A4(n338), .ZN(
        decodeReadData1_o[45]) );
  CKND2D0 U1111 ( .A1(n1099), .A2(\completionDataOut[4][39] ), .ZN(n547) );
  CKND2D0 U1112 ( .A1(n1116), .A2(\completionDataOut[6][39] ), .ZN(n548) );
  CKND2D0 U1113 ( .A1(n1099), .A2(\completionDataOut[4][38] ), .ZN(n550) );
  CKND2D0 U1114 ( .A1(n1116), .A2(\completionDataOut[6][38] ), .ZN(n551) );
  CKND2D0 U1115 ( .A1(n1100), .A2(\completionDataOut[4][30] ), .ZN(n553) );
  CKND2D0 U1116 ( .A1(n1111), .A2(\completionDataOut[6][30] ), .ZN(n554) );
  CKND2D0 U1117 ( .A1(n1107), .A2(\completionDataOut[4][28] ), .ZN(n556) );
  CKND2D0 U1118 ( .A1(n1112), .A2(\completionDataOut[6][28] ), .ZN(n557) );
  CKND2D0 U1119 ( .A1(n1105), .A2(\completionDataOut[4][25] ), .ZN(n559) );
  CKND2D0 U1120 ( .A1(n1112), .A2(\completionDataOut[6][25] ), .ZN(n560) );
  CKND2D0 U1121 ( .A1(n1104), .A2(\completionDataOut[4][13] ), .ZN(n562) );
  CKND2D0 U1122 ( .A1(n1119), .A2(\completionDataOut[6][13] ), .ZN(n563) );
  CKND2D0 U1123 ( .A1(n1103), .A2(\completionDataOut[4][9] ), .ZN(n565) );
  CKND2D0 U1124 ( .A1(n1114), .A2(\completionDataOut[6][9] ), .ZN(n566) );
  CKND2D0 U1125 ( .A1(n1102), .A2(\completionDataOut[4][5] ), .ZN(n568) );
  CKND2D0 U1126 ( .A1(n1114), .A2(\completionDataOut[6][5] ), .ZN(n569) );
  CKND2D0 U1127 ( .A1(n1102), .A2(\completionDataOut[4][4] ), .ZN(n571) );
  CKND2D0 U1128 ( .A1(n1115), .A2(\completionDataOut[6][4] ), .ZN(n572) );
  CKND2D0 U1129 ( .A1(n1207), .A2(\completionDataOut[4][59] ), .ZN(n574) );
  CKND2D0 U1130 ( .A1(n1209), .A2(\completionDataOut[6][59] ), .ZN(n575) );
  CKND2D0 U1131 ( .A1(n1197), .A2(\completionDataOut[4][53] ), .ZN(n577) );
  CKND2D0 U1132 ( .A1(n1210), .A2(\completionDataOut[6][53] ), .ZN(n578) );
  CKND2D0 U1133 ( .A1(n1198), .A2(\completionDataOut[4][50] ), .ZN(n580) );
  CKND2D0 U1134 ( .A1(n1218), .A2(\completionDataOut[6][50] ), .ZN(n581) );
  CKND2D0 U1135 ( .A1(n1198), .A2(\completionDataOut[4][47] ), .ZN(n583) );
  CKND2D0 U1136 ( .A1(n1219), .A2(\completionDataOut[6][47] ), .ZN(n584) );
  CKND2D0 U1137 ( .A1(n1199), .A2(\completionDataOut[4][41] ), .ZN(n586) );
  CKND2D0 U1138 ( .A1(n1211), .A2(\completionDataOut[6][41] ), .ZN(n587) );
  CKND2D0 U1139 ( .A1(n1200), .A2(\completionDataOut[4][37] ), .ZN(n589) );
  CKND2D0 U1140 ( .A1(n1217), .A2(\completionDataOut[6][37] ), .ZN(n590) );
  CKND2D0 U1141 ( .A1(n1200), .A2(\completionDataOut[4][35] ), .ZN(n592) );
  CKND2D0 U1142 ( .A1(n1217), .A2(\completionDataOut[6][35] ), .ZN(n593) );
  CKND2D0 U1143 ( .A1(n1201), .A2(\completionDataOut[4][29] ), .ZN(n595) );
  CKND2D0 U1144 ( .A1(n1212), .A2(\completionDataOut[6][29] ), .ZN(n596) );
  CKND2D0 U1145 ( .A1(n1206), .A2(\completionDataOut[4][23] ), .ZN(n598) );
  CKND2D0 U1146 ( .A1(n1213), .A2(\completionDataOut[6][23] ), .ZN(n599) );
  CKND2D0 U1147 ( .A1(n1202), .A2(\completionDataOut[4][17] ), .ZN(n601) );
  CKND2D0 U1148 ( .A1(n1214), .A2(\completionDataOut[6][17] ), .ZN(n602) );
  CKND2D0 U1149 ( .A1(n1208), .A2(\completionDataOut[4][15] ), .ZN(n604) );
  CKND2D0 U1150 ( .A1(n1221), .A2(\completionDataOut[6][15] ), .ZN(n605) );
  CKND2D0 U1151 ( .A1(n1205), .A2(\completionDataOut[4][11] ), .ZN(n607) );
  CKND2D0 U1152 ( .A1(n1220), .A2(\completionDataOut[6][11] ), .ZN(n608) );
  CKND2D0 U1153 ( .A1(n1204), .A2(\completionDataOut[4][8] ), .ZN(n610) );
  CKND2D0 U1154 ( .A1(n1215), .A2(\completionDataOut[6][8] ), .ZN(n611) );
  CKND2D0 U1155 ( .A1(n1203), .A2(\completionDataOut[4][3] ), .ZN(n613) );
  CKND2D0 U1156 ( .A1(n1216), .A2(\completionDataOut[6][3] ), .ZN(n614) );
  CKND2D0 U1157 ( .A1(n1203), .A2(\completionDataOut[4][2] ), .ZN(n616) );
  CKND2D0 U1158 ( .A1(n1216), .A2(\completionDataOut[6][2] ), .ZN(n617) );
  CKND2D0 U1159 ( .A1(n986), .A2(\completionDataOut[4][61] ), .ZN(n619) );
  CKND2D0 U1160 ( .A1(n1003), .A2(\completionDataOut[6][61] ), .ZN(n620) );
  CKND2D0 U1161 ( .A1(n986), .A2(\completionDataOut[4][60] ), .ZN(n622) );
  CKND2D0 U1162 ( .A1(n1003), .A2(\completionDataOut[6][60] ), .ZN(n623) );
  CKND2D0 U1163 ( .A1(n989), .A2(\completionDataOut[4][56] ), .ZN(n625) );
  CKND2D0 U1164 ( .A1(n1006), .A2(\completionDataOut[6][56] ), .ZN(n626) );
  ND4D8 U1165 ( .A1(n1396), .A2(n528), .A3(n624), .A4(n337), .ZN(
        commitReadData_o[56]) );
  CKND2D0 U1166 ( .A1(n989), .A2(\completionDataOut[4][55] ), .ZN(n628) );
  CKND2D0 U1167 ( .A1(n1008), .A2(\completionDataOut[6][55] ), .ZN(n629) );
  CKND2D0 U1168 ( .A1(n985), .A2(\completionDataOut[4][49] ), .ZN(n631) );
  CKND2D0 U1169 ( .A1(n1002), .A2(\completionDataOut[6][49] ), .ZN(n632) );
  CKND2D0 U1170 ( .A1(n985), .A2(\completionDataOut[4][48] ), .ZN(n634) );
  CKND2D0 U1171 ( .A1(n1002), .A2(\completionDataOut[6][48] ), .ZN(n635) );
  CKND2D0 U1172 ( .A1(n990), .A2(\completionDataOut[4][44] ), .ZN(n637) );
  CKND2D0 U1173 ( .A1(n1011), .A2(\completionDataOut[6][44] ), .ZN(n638) );
  ND4D8 U1174 ( .A1(n1435), .A2(n1436), .A3(n636), .A4(n334), .ZN(
        commitReadData_o[44]) );
  CKND2D0 U1175 ( .A1(n990), .A2(\completionDataOut[4][43] ), .ZN(n640) );
  CKND2D0 U1176 ( .A1(n1007), .A2(\completionDataOut[6][43] ), .ZN(n641) );
  CKND2D0 U1177 ( .A1(n984), .A2(\completionDataOut[4][36] ), .ZN(n643) );
  CKND2D0 U1178 ( .A1(n1001), .A2(\completionDataOut[6][36] ), .ZN(n644) );
  CKND2D0 U1179 ( .A1(n991), .A2(\completionDataOut[4][31] ), .ZN(n646) );
  CKND2D0 U1180 ( .A1(n1000), .A2(\completionDataOut[6][31] ), .ZN(n647) );
  CKND2D0 U1181 ( .A1(n983), .A2(\completionDataOut[4][24] ), .ZN(n649) );
  CKND2D0 U1182 ( .A1(n999), .A2(\completionDataOut[6][24] ), .ZN(n650) );
  CKND2D0 U1183 ( .A1(n995), .A2(\completionDataOut[4][19] ), .ZN(n652) );
  CKND2D0 U1184 ( .A1(n1009), .A2(\completionDataOut[6][19] ), .ZN(n653) );
  CKND2D0 U1185 ( .A1(n993), .A2(\completionDataOut[4][18] ), .ZN(n655) );
  CKND2D0 U1186 ( .A1(n1012), .A2(\completionDataOut[6][18] ), .ZN(n656) );
  CKND2D0 U1187 ( .A1(n982), .A2(\completionDataOut[4][12] ), .ZN(n658) );
  CKND2D0 U1188 ( .A1(n998), .A2(\completionDataOut[6][12] ), .ZN(n659) );
  CKND2D0 U1189 ( .A1(n992), .A2(\completionDataOut[4][7] ), .ZN(n661) );
  CKND2D0 U1190 ( .A1(n1010), .A2(\completionDataOut[6][7] ), .ZN(n662) );
  CKND2D0 U1191 ( .A1(n981), .A2(\completionDataOut[4][1] ), .ZN(n664) );
  CKND2D0 U1192 ( .A1(n997), .A2(\completionDataOut[6][1] ), .ZN(n665) );
  CKND2D0 U1193 ( .A1(n981), .A2(\completionDataOut[4][0] ), .ZN(n667) );
  CKND2D0 U1194 ( .A1(n997), .A2(\completionDataOut[6][0] ), .ZN(n668) );
  CKND2D0 U1195 ( .A1(n1130), .A2(\completionDataOut[5][62] ), .ZN(n670) );
  CKND2D0 U1196 ( .A1(n1133), .A2(\completionDataOut[7][62] ), .ZN(n671) );
  CKND2D0 U1197 ( .A1(n1120), .A2(\completionDataOut[5][54] ), .ZN(n673) );
  CKND2D0 U1198 ( .A1(n1134), .A2(\completionDataOut[7][54] ), .ZN(n674) );
  ND4D8 U1199 ( .A1(n1786), .A2(n130), .A3(n534), .A4(n672), .ZN(
        decodeReadData1_o[54]) );
  CKND2D0 U1200 ( .A1(n1121), .A2(\completionDataOut[5][52] ), .ZN(n676) );
  CKND2D0 U1201 ( .A1(n1143), .A2(\completionDataOut[7][52] ), .ZN(n677) );
  ND4D8 U1202 ( .A1(n1780), .A2(n131), .A3(n537), .A4(n675), .ZN(
        decodeReadData1_o[52]) );
  CKND2D0 U1203 ( .A1(n1121), .A2(\completionDataOut[5][51] ), .ZN(n679) );
  CKND2D0 U1204 ( .A1(n1142), .A2(\completionDataOut[7][51] ), .ZN(n680) );
  ND4D8 U1205 ( .A1(n1779), .A2(n25), .A3(n540), .A4(n678), .ZN(
        decodeReadData1_o[51]) );
  CKND2D0 U1206 ( .A1(n1122), .A2(\completionDataOut[5][44] ), .ZN(n682) );
  CKND2D0 U1207 ( .A1(n1135), .A2(\completionDataOut[7][44] ), .ZN(n683) );
  CKND2D0 U1208 ( .A1(n1123), .A2(\completionDataOut[5][39] ), .ZN(n685) );
  CKND2D0 U1209 ( .A1(n1141), .A2(\completionDataOut[7][39] ), .ZN(n686) );
  ND4D8 U1210 ( .A1(n1737), .A2(n137), .A3(n546), .A4(n684), .ZN(
        decodeReadData1_o[39]) );
  CKND2D0 U1211 ( .A1(n1123), .A2(\completionDataOut[5][38] ), .ZN(n688) );
  CKND2D0 U1212 ( .A1(n1141), .A2(\completionDataOut[7][38] ), .ZN(n689) );
  ND4D8 U1213 ( .A1(n1736), .A2(n26), .A3(n549), .A4(n687), .ZN(
        decodeReadData1_o[38]) );
  CKND2D0 U1214 ( .A1(n1124), .A2(\completionDataOut[5][30] ), .ZN(n691) );
  CKND2D0 U1215 ( .A1(n1136), .A2(\completionDataOut[7][30] ), .ZN(n692) );
  ND4D8 U1216 ( .A1(n1706), .A2(n140), .A3(n552), .A4(n690), .ZN(
        decodeReadData1_o[30]) );
  CKND2D0 U1217 ( .A1(n1131), .A2(\completionDataOut[5][28] ), .ZN(n694) );
  CKND2D0 U1218 ( .A1(n1137), .A2(\completionDataOut[7][28] ), .ZN(n695) );
  ND4D8 U1219 ( .A1(n1700), .A2(n141), .A3(n555), .A4(n693), .ZN(
        decodeReadData1_o[28]) );
  CKND2D0 U1220 ( .A1(n1129), .A2(\completionDataOut[5][25] ), .ZN(n697) );
  CKND2D0 U1221 ( .A1(n1137), .A2(\completionDataOut[7][25] ), .ZN(n698) );
  ND4D8 U1222 ( .A1(n1691), .A2(n27), .A3(n558), .A4(n696), .ZN(
        decodeReadData1_o[25]) );
  CKND2D0 U1223 ( .A1(n1125), .A2(\completionDataOut[5][18] ), .ZN(n700) );
  CKND2D0 U1224 ( .A1(n1138), .A2(\completionDataOut[7][18] ), .ZN(n701) );
  ND4D8 U1225 ( .A1(n1665), .A2(n513), .A3(n170), .A4(n699), .ZN(
        decodeReadData1_o[18]) );
  CKND2D0 U1226 ( .A1(n1128), .A2(\completionDataOut[5][13] ), .ZN(n703) );
  CKND2D0 U1227 ( .A1(n1144), .A2(\completionDataOut[7][13] ), .ZN(n704) );
  ND4D8 U1228 ( .A1(n1648), .A2(n28), .A3(n561), .A4(n702), .ZN(
        decodeReadData1_o[13]) );
  CKND2D0 U1229 ( .A1(n1127), .A2(\completionDataOut[5][9] ), .ZN(n706) );
  CKND2D0 U1230 ( .A1(n1139), .A2(\completionDataOut[7][9] ), .ZN(n707) );
  ND4D8 U1231 ( .A1(n1634), .A2(n146), .A3(n564), .A4(n705), .ZN(
        decodeReadData1_o[9]) );
  CKND2D0 U1232 ( .A1(n1126), .A2(\completionDataOut[5][5] ), .ZN(n709) );
  CKND2D0 U1233 ( .A1(n1139), .A2(\completionDataOut[7][5] ), .ZN(n710) );
  ND4D8 U1234 ( .A1(n1621), .A2(n29), .A3(n567), .A4(n708), .ZN(
        decodeReadData1_o[5]) );
  CKND2D0 U1235 ( .A1(n1126), .A2(\completionDataOut[5][4] ), .ZN(n712) );
  CKND2D0 U1236 ( .A1(n1140), .A2(\completionDataOut[7][4] ), .ZN(n713) );
  ND4D8 U1237 ( .A1(n1620), .A2(n31), .A3(n570), .A4(n711), .ZN(
        decodeReadData1_o[4]) );
  CKND2D0 U1238 ( .A1(n1232), .A2(\completionDataOut[5][59] ), .ZN(n715) );
  CKND2D0 U1239 ( .A1(n1234), .A2(\completionDataOut[7][59] ), .ZN(n716) );
  ND4D8 U1240 ( .A1(n2039), .A2(n151), .A3(n573), .A4(n714), .ZN(
        decodeReadData2_o[59]) );
  CKND2D0 U1241 ( .A1(n1222), .A2(\completionDataOut[5][53] ), .ZN(n718) );
  CKND2D0 U1242 ( .A1(n1235), .A2(\completionDataOut[7][53] ), .ZN(n719) );
  ND4D8 U1243 ( .A1(n2017), .A2(n152), .A3(n576), .A4(n717), .ZN(
        decodeReadData2_o[53]) );
  CKND2D0 U1244 ( .A1(n1223), .A2(\completionDataOut[5][50] ), .ZN(n721) );
  CKND2D0 U1245 ( .A1(n1243), .A2(\completionDataOut[7][50] ), .ZN(n722) );
  ND4D8 U1246 ( .A1(n2007), .A2(n153), .A3(n579), .A4(n720), .ZN(
        decodeReadData2_o[50]) );
  CKND2D0 U1247 ( .A1(n1223), .A2(\completionDataOut[5][47] ), .ZN(n724) );
  CKND2D0 U1248 ( .A1(n1244), .A2(\completionDataOut[7][47] ), .ZN(n725) );
  ND4D8 U1249 ( .A1(n1998), .A2(n32), .A3(n582), .A4(n723), .ZN(
        decodeReadData2_o[47]) );
  CKND2D0 U1250 ( .A1(n1224), .A2(\completionDataOut[5][41] ), .ZN(n727) );
  CKND2D0 U1251 ( .A1(n1236), .A2(\completionDataOut[7][41] ), .ZN(n728) );
  ND4D8 U1252 ( .A1(n1976), .A2(n156), .A3(n585), .A4(n726), .ZN(
        decodeReadData2_o[41]) );
  CKND2D0 U1253 ( .A1(n1225), .A2(\completionDataOut[5][37] ), .ZN(n730) );
  CKND2D0 U1254 ( .A1(n1242), .A2(\completionDataOut[7][37] ), .ZN(n731) );
  ND4D8 U1255 ( .A1(n1962), .A2(n1963), .A3(n588), .A4(n729), .ZN(
        decodeReadData2_o[37]) );
  CKND2D0 U1256 ( .A1(n1225), .A2(\completionDataOut[5][35] ), .ZN(n733) );
  CKND2D0 U1257 ( .A1(n1242), .A2(\completionDataOut[7][35] ), .ZN(n734) );
  ND4D8 U1258 ( .A1(n1956), .A2(n1957), .A3(n591), .A4(n732), .ZN(
        decodeReadData2_o[35]) );
  CKND2D0 U1259 ( .A1(n1226), .A2(\completionDataOut[5][29] ), .ZN(n736) );
  CKND2D0 U1260 ( .A1(n1237), .A2(\completionDataOut[7][29] ), .ZN(n737) );
  ND4D8 U1261 ( .A1(n1935), .A2(n33), .A3(n594), .A4(n735), .ZN(
        decodeReadData2_o[29]) );
  CKND2D0 U1262 ( .A1(n1231), .A2(\completionDataOut[5][23] ), .ZN(n739) );
  CKND2D0 U1263 ( .A1(n1238), .A2(\completionDataOut[7][23] ), .ZN(n740) );
  ND4D8 U1264 ( .A1(n1914), .A2(n34), .A3(n597), .A4(n738), .ZN(
        decodeReadData2_o[23]) );
  CKND2D0 U1265 ( .A1(n1227), .A2(\completionDataOut[5][17] ), .ZN(n742) );
  CKND2D0 U1266 ( .A1(n1239), .A2(\completionDataOut[7][17] ), .ZN(n743) );
  ND4D8 U1267 ( .A1(n1892), .A2(n100), .A3(n600), .A4(n741), .ZN(
        decodeReadData2_o[17]) );
  CKND2D0 U1268 ( .A1(n1233), .A2(\completionDataOut[5][15] ), .ZN(n745) );
  CKND2D0 U1269 ( .A1(n1246), .A2(\completionDataOut[7][15] ), .ZN(n746) );
  ND4D8 U1270 ( .A1(n1886), .A2(n101), .A3(n603), .A4(n744), .ZN(
        decodeReadData2_o[15]) );
  CKND2D0 U1271 ( .A1(n1230), .A2(\completionDataOut[5][11] ), .ZN(n748) );
  CKND2D0 U1272 ( .A1(n1245), .A2(\completionDataOut[7][11] ), .ZN(n749) );
  ND4D8 U1273 ( .A1(n1872), .A2(n102), .A3(n606), .A4(n747), .ZN(
        decodeReadData2_o[11]) );
  CKND2D0 U1274 ( .A1(n1229), .A2(\completionDataOut[5][8] ), .ZN(n751) );
  CKND2D0 U1275 ( .A1(n1240), .A2(\completionDataOut[7][8] ), .ZN(n752) );
  ND4D8 U1276 ( .A1(n1863), .A2(n35), .A3(n609), .A4(n750), .ZN(
        decodeReadData2_o[8]) );
  CKND2D0 U1277 ( .A1(n1228), .A2(\completionDataOut[5][3] ), .ZN(n754) );
  CKND2D0 U1278 ( .A1(n1241), .A2(\completionDataOut[7][3] ), .ZN(n755) );
  ND4D8 U1279 ( .A1(n1845), .A2(n105), .A3(n612), .A4(n753), .ZN(
        decodeReadData2_o[3]) );
  CKND2D0 U1280 ( .A1(n1228), .A2(\completionDataOut[5][2] ), .ZN(n757) );
  CKND2D0 U1281 ( .A1(n1241), .A2(\completionDataOut[7][2] ), .ZN(n758) );
  ND4D8 U1282 ( .A1(n1844), .A2(n36), .A3(n615), .A4(n756), .ZN(
        decodeReadData2_o[2]) );
  CKND2D0 U1283 ( .A1(n1018), .A2(\completionDataOut[5][61] ), .ZN(n760) );
  CKND2D0 U1284 ( .A1(n1035), .A2(\completionDataOut[7][61] ), .ZN(n761) );
  ND4D8 U1285 ( .A1(n1382), .A2(n97), .A3(n618), .A4(n759), .ZN(
        commitReadData_o[61]) );
  CKND2D0 U1286 ( .A1(n1018), .A2(\completionDataOut[5][60] ), .ZN(n763) );
  CKND2D0 U1287 ( .A1(n1035), .A2(\completionDataOut[7][60] ), .ZN(n764) );
  ND4D8 U1288 ( .A1(n1384), .A2(n98), .A3(n621), .A4(n762), .ZN(
        commitReadData_o[60]) );
  CKND2D0 U1289 ( .A1(n1021), .A2(\completionDataOut[5][55] ), .ZN(n766) );
  CKND2D0 U1290 ( .A1(n1040), .A2(\completionDataOut[7][55] ), .ZN(n767) );
  ND4D8 U1291 ( .A1(n1398), .A2(n108), .A3(n627), .A4(n765), .ZN(
        commitReadData_o[55]) );
  CKND2D0 U1292 ( .A1(n1017), .A2(\completionDataOut[5][49] ), .ZN(n769) );
  CKND2D0 U1293 ( .A1(n1034), .A2(\completionDataOut[7][49] ), .ZN(n770) );
  ND4D8 U1294 ( .A1(n1420), .A2(n109), .A3(n630), .A4(n768), .ZN(
        commitReadData_o[49]) );
  CKND2D0 U1295 ( .A1(n1017), .A2(\completionDataOut[5][48] ), .ZN(n772) );
  CKND2D0 U1296 ( .A1(n1034), .A2(\completionDataOut[7][48] ), .ZN(n773) );
  ND4D8 U1297 ( .A1(n1422), .A2(n110), .A3(n633), .A4(n771), .ZN(
        commitReadData_o[48]) );
  CKND2D0 U1298 ( .A1(n1022), .A2(\completionDataOut[5][43] ), .ZN(n775) );
  CKND2D0 U1299 ( .A1(n1039), .A2(\completionDataOut[7][43] ), .ZN(n776) );
  ND4D8 U1300 ( .A1(n1438), .A2(n37), .A3(n639), .A4(n774), .ZN(
        commitReadData_o[43]) );
  CKND2D0 U1301 ( .A1(n1026), .A2(\completionDataOut[5][42] ), .ZN(n778) );
  CKND2D0 U1302 ( .A1(n1043), .A2(\completionDataOut[7][42] ), .ZN(n779) );
  CKND2D0 U1303 ( .A1(n1016), .A2(\completionDataOut[5][36] ), .ZN(n781) );
  CKND2D0 U1304 ( .A1(n1033), .A2(\completionDataOut[7][36] ), .ZN(n782) );
  ND4D8 U1305 ( .A1(n1462), .A2(n113), .A3(n642), .A4(n780), .ZN(
        commitReadData_o[36]) );
  CKND2D0 U1306 ( .A1(n1023), .A2(\completionDataOut[5][31] ), .ZN(n784) );
  CKND2D0 U1307 ( .A1(n1032), .A2(\completionDataOut[7][31] ), .ZN(n785) );
  ND4D8 U1308 ( .A1(n1480), .A2(n1481), .A3(n645), .A4(n783), .ZN(
        commitReadData_o[31]) );
  CKND2D0 U1309 ( .A1(n1015), .A2(\completionDataOut[5][24] ), .ZN(n787) );
  CKND2D0 U1310 ( .A1(n1031), .A2(\completionDataOut[7][24] ), .ZN(n788) );
  ND4D8 U1311 ( .A1(n1506), .A2(n118), .A3(n648), .A4(n786), .ZN(
        commitReadData_o[24]) );
  CKND2D0 U1312 ( .A1(n1027), .A2(\completionDataOut[5][19] ), .ZN(n790) );
  CKND2D0 U1313 ( .A1(n1041), .A2(\completionDataOut[7][19] ), .ZN(n791) );
  ND4D8 U1314 ( .A1(n1524), .A2(n38), .A3(n651), .A4(n789), .ZN(
        commitReadData_o[19]) );
  CKND2D0 U1315 ( .A1(n1014), .A2(\completionDataOut[5][12] ), .ZN(n793) );
  CKND2D0 U1316 ( .A1(n1030), .A2(\completionDataOut[7][12] ), .ZN(n794) );
  ND4D8 U1317 ( .A1(n1548), .A2(n1549), .A3(n657), .A4(n792), .ZN(
        commitReadData_o[12]) );
  CKND2D0 U1318 ( .A1(n1024), .A2(\completionDataOut[5][7] ), .ZN(n796) );
  CKND2D0 U1319 ( .A1(n1042), .A2(\completionDataOut[7][7] ), .ZN(n797) );
  ND4D8 U1320 ( .A1(n1566), .A2(n39), .A3(n660), .A4(n795), .ZN(
        commitReadData_o[7]) );
  CKND2D0 U1321 ( .A1(n1025), .A2(\completionDataOut[5][6] ), .ZN(n799) );
  CKND2D0 U1322 ( .A1(n1044), .A2(\completionDataOut[7][6] ), .ZN(n800) );
  CKND2D0 U1323 ( .A1(n1013), .A2(\completionDataOut[5][1] ), .ZN(n802) );
  CKND2D0 U1324 ( .A1(n1029), .A2(\completionDataOut[7][1] ), .ZN(n803) );
  ND4D8 U1325 ( .A1(n1586), .A2(n128), .A3(n663), .A4(n801), .ZN(
        commitReadData_o[1]) );
  CKND2D0 U1326 ( .A1(n1013), .A2(\completionDataOut[5][0] ), .ZN(n805) );
  CKND2D0 U1327 ( .A1(n1029), .A2(\completionDataOut[7][0] ), .ZN(n806) );
  ND4D8 U1328 ( .A1(n1588), .A2(n129), .A3(n666), .A4(n804), .ZN(
        commitReadData_o[0]) );
  ND4D8 U1329 ( .A1(n1332), .A2(n1333), .A3(n1334), .A4(n324), .ZN(
        commitReadData_o[74]) );
  ND4D8 U1330 ( .A1(n1340), .A2(n1341), .A3(n1342), .A4(n1343), .ZN(
        commitReadData_o[72]) );
  AOI22D2 U1331 ( .A1(n1028), .A2(\managementDataOut[5][2] ), .B1(n1040), .B2(
        \managementDataOut[7][2] ), .ZN(n1343) );
  ND4D8 U1332 ( .A1(n1348), .A2(n1349), .A3(n1350), .A4(n325), .ZN(
        commitReadData_o[70]) );
  ND4D8 U1333 ( .A1(n1352), .A2(n1353), .A3(n1354), .A4(n326), .ZN(
        commitReadData_o[69]) );
  ND4D8 U1334 ( .A1(n1356), .A2(n1357), .A3(n1358), .A4(n327), .ZN(
        commitReadData_o[68]) );
  ND4D8 U1335 ( .A1(n1360), .A2(n1361), .A3(n1362), .A4(n328), .ZN(
        commitReadData_o[67]) );
  ND4D8 U1336 ( .A1(n1364), .A2(n1365), .A3(n1366), .A4(n329), .ZN(
        commitReadData_o[66]) );
  ND4D8 U1337 ( .A1(n1368), .A2(n1369), .A3(n1370), .A4(n1371), .ZN(
        commitReadData_o[65]) );
  CKND2D0 U1338 ( .A1(commitReadAddr_i[0]), .A2(commitReadAddr_i[1]), .ZN(
        n1310) );
  CKND2D0 U1339 ( .A1(commitReadAddr_i[0]), .A2(n1591), .ZN(n1308) );
  CKND0 U1340 ( .I(commitReadAddr_i[1]), .ZN(n1591) );
  CKND2D0 U1341 ( .A1(commitReadAddr_i[1]), .A2(n1590), .ZN(n1306) );
  CKND0 U1342 ( .I(commitReadAddr_i[0]), .ZN(n1590) );
  AO22D0 U1343 ( .A1(n221), .A2(n916), .B1(n1275), .B2(
        \completionDataOut[6][26] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[26].enDff/theFlop/N3 )
         );
  AO22D0 U1344 ( .A1(completionWriteData_i[20]), .A2(n942), .B1(n928), .B2(
        \completionDataOut[7][20] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[20].enDff/theFlop/N3 )
         );
  AO22D0 U1345 ( .A1(n199), .A2(n912), .B1(n903), .B2(
        \completionDataOut[6][4] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U1346 ( .A1(n245), .A2(n912), .B1(n903), .B2(
        \completionDataOut[6][50] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[50].enDff/theFlop/N3 )
         );
  CKBD1 U1347 ( .I(n192), .Z(n1248) );
  AO22D0 U1348 ( .A1(n834), .A2(\completionDataOut[2][48] ), .B1(n811), .B2(
        completionWriteData_i[48]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[48].enDff/theFlop/N3 )
         );
  AO22D0 U1349 ( .A1(completionWriteData_i[26]), .A2(n889), .B1(n875), .B2(
        \completionDataOut[5][26] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[26].enDff/theFlop/N3 )
         );
  AO22D0 U1350 ( .A1(n830), .A2(\completionDataOut[2][41] ), .B1(n812), .B2(
        completionWriteData_i[41]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[41].enDff/theFlop/N3 )
         );
  AO22D0 U1351 ( .A1(n830), .A2(\completionDataOut[2][40] ), .B1(n812), .B2(
        completionWriteData_i[40]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[40].enDff/theFlop/N3 )
         );
  AO22D0 U1352 ( .A1(n827), .A2(\completionDataOut[2][67] ), .B1(n821), .B2(
        completionWriteData_i[67]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[67].enDff/theFlop/N3 )
         );
  AO22D0 U1353 ( .A1(n215), .A2(n862), .B1(n847), .B2(
        \completionDataOut[3][20] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[20].enDff/theFlop/N3 )
         );
  AO22D0 U1354 ( .A1(n210), .A2(n916), .B1(n900), .B2(
        \completionDataOut[6][15] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[15].enDff/theFlop/N3 )
         );
  AO22D0 U1355 ( .A1(n224), .A2(n914), .B1(n902), .B2(
        \completionDataOut[6][29] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[29].enDff/theFlop/N3 )
         );
  AO22D0 U1356 ( .A1(n222), .A2(n914), .B1(n1275), .B2(
        \completionDataOut[6][27] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[27].enDff/theFlop/N3 )
         );
  AO22D0 U1357 ( .A1(n223), .A2(n914), .B1(n902), .B2(
        \completionDataOut[6][28] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[28].enDff/theFlop/N3 )
         );
  AO22D0 U1358 ( .A1(n212), .A2(n915), .B1(n898), .B2(
        \completionDataOut[6][17] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[17].enDff/theFlop/N3 )
         );
  AO22D0 U1359 ( .A1(completionWriteData_i[16]), .A2(n915), .B1(n903), .B2(
        \completionDataOut[6][16] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[16].enDff/theFlop/N3 )
         );
  AO22D0 U1360 ( .A1(n213), .A2(n915), .B1(n1275), .B2(
        \completionDataOut[6][18] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[18].enDff/theFlop/N3 )
         );
  AO22D0 U1361 ( .A1(n214), .A2(n915), .B1(n901), .B2(
        \completionDataOut[6][19] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[19].enDff/theFlop/N3 )
         );
  AO22D0 U1362 ( .A1(n196), .A2(n915), .B1(n899), .B2(
        \completionDataOut[6][1] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U1363 ( .A1(n831), .A2(\completionDataOut[2][29] ), .B1(n820), .B2(
        completionWriteData_i[29]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[29].enDff/theFlop/N3 )
         );
  AO22D0 U1364 ( .A1(n830), .A2(\completionDataOut[2][3] ), .B1(n820), .B2(
        completionWriteData_i[3]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U1365 ( .A1(n827), .A2(\completionDataOut[2][66] ), .B1(n820), .B2(
        completionWriteData_i[66]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[66].enDff/theFlop/N3 )
         );
  AO22D0 U1366 ( .A1(completionWriteData_i[21]), .A2(n940), .B1(n928), .B2(
        \completionDataOut[7][21] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[21].enDff/theFlop/N3 )
         );
  AO22D0 U1367 ( .A1(n245), .A2(n933), .B1(n929), .B2(
        \completionDataOut[7][50] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[50].enDff/theFlop/N3 )
         );
  AO22D0 U1368 ( .A1(n199), .A2(n933), .B1(n929), .B2(
        \completionDataOut[7][4] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U1369 ( .A1(completionWriteData_i[15]), .A2(n889), .B1(n864), .B2(
        \completionDataOut[5][15] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[15].enDff/theFlop/N3 )
         );
  AO22D0 U1370 ( .A1(n225), .A2(n914), .B1(n899), .B2(
        \completionDataOut[6][30] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[30].enDff/theFlop/N3 )
         );
  AO22D0 U1371 ( .A1(n197), .A2(n914), .B1(n901), .B2(
        \completionDataOut[6][2] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U1372 ( .A1(completionWriteData_i[27]), .A2(n887), .B1(n875), .B2(
        \completionDataOut[5][27] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[27].enDff/theFlop/N3 )
         );
  AO22D0 U1373 ( .A1(completionWriteData_i[1]), .A2(n888), .B1(n864), .B2(
        \completionDataOut[5][1] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U1374 ( .A1(completionWriteData_i[19]), .A2(n888), .B1(n864), .B2(
        \completionDataOut[5][19] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[19].enDff/theFlop/N3 )
         );
  AO22D0 U1375 ( .A1(completionWriteData_i[18]), .A2(n888), .B1(n864), .B2(
        \completionDataOut[5][18] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[18].enDff/theFlop/N3 )
         );
  AO22D0 U1376 ( .A1(n211), .A2(n888), .B1(n864), .B2(
        \completionDataOut[5][16] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[16].enDff/theFlop/N3 )
         );
  AO22D0 U1377 ( .A1(completionWriteData_i[29]), .A2(n887), .B1(n875), .B2(
        \completionDataOut[5][29] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[29].enDff/theFlop/N3 )
         );
  AO22D0 U1378 ( .A1(completionWriteData_i[17]), .A2(n888), .B1(n864), .B2(
        \completionDataOut[5][17] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[17].enDff/theFlop/N3 )
         );
  AO22D0 U1379 ( .A1(completionWriteData_i[28]), .A2(n887), .B1(n875), .B2(
        \completionDataOut[5][28] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[28].enDff/theFlop/N3 )
         );
  AO22D0 U1380 ( .A1(completionWriteData_i[45]), .A2(n880), .B1(n876), .B2(
        \completionDataOut[5][45] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[45].enDff/theFlop/N3 )
         );
  AO22D0 U1381 ( .A1(completionWriteData_i[44]), .A2(n880), .B1(n876), .B2(
        \completionDataOut[5][44] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[44].enDff/theFlop/N3 )
         );
  AO22D0 U1382 ( .A1(n827), .A2(\completionDataOut[2][64] ), .B1(n819), .B2(
        completionWriteData_i[64]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[64].enDff/theFlop/N3 )
         );
  AO22D0 U1383 ( .A1(n829), .A2(\completionDataOut[2][4] ), .B1(n811), .B2(
        completionWriteData_i[4]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U1384 ( .A1(n829), .A2(\completionDataOut[2][50] ), .B1(n811), .B2(
        completionWriteData_i[50]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[50].enDff/theFlop/N3 )
         );
  AO22D0 U1385 ( .A1(n828), .A2(\completionDataOut[2][63] ), .B1(n819), .B2(
        completionWriteData_i[63]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[63].enDff/theFlop/N3 )
         );
  AO22D0 U1386 ( .A1(n828), .A2(\completionDataOut[2][62] ), .B1(n819), .B2(
        completionWriteData_i[62]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[62].enDff/theFlop/N3 )
         );
  AO22D0 U1387 ( .A1(n829), .A2(\completionDataOut[2][49] ), .B1(n811), .B2(
        completionWriteData_i[49]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[49].enDff/theFlop/N3 )
         );
  AO22D0 U1388 ( .A1(n201), .A2(n910), .B1(n898), .B2(
        \completionDataOut[6][6] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U1389 ( .A1(n244), .A2(n912), .B1(n900), .B2(
        \completionDataOut[6][49] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[49].enDff/theFlop/N3 )
         );
  AO22D0 U1390 ( .A1(n246), .A2(n912), .B1(n900), .B2(
        \completionDataOut[6][51] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[51].enDff/theFlop/N3 )
         );
  AO22D0 U1391 ( .A1(n203), .A2(n910), .B1(n898), .B2(
        \completionDataOut[6][8] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U1392 ( .A1(n247), .A2(n912), .B1(n900), .B2(
        \completionDataOut[6][52] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[52].enDff/theFlop/N3 )
         );
  AO22D0 U1393 ( .A1(n202), .A2(n910), .B1(n898), .B2(
        \completionDataOut[6][7] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U1394 ( .A1(n204), .A2(n910), .B1(n898), .B2(
        \completionDataOut[6][9] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[9].enDff/theFlop/N3 ) );
  AO22D0 U1395 ( .A1(n207), .A2(n941), .B1(n924), .B2(
        \completionDataOut[7][12] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[12].enDff/theFlop/N3 )
         );
  AO22D0 U1396 ( .A1(n208), .A2(n941), .B1(n929), .B2(
        \completionDataOut[7][13] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[13].enDff/theFlop/N3 )
         );
  AO22D0 U1397 ( .A1(n195), .A2(n942), .B1(n926), .B2(
        \completionDataOut[7][0] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U1398 ( .A1(completionWriteData_i[10]), .A2(n941), .B1(n927), .B2(
        \completionDataOut[7][10] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[10].enDff/theFlop/N3 )
         );
  AO22D0 U1399 ( .A1(n209), .A2(n941), .B1(n925), .B2(
        \completionDataOut[7][14] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[14].enDff/theFlop/N3 )
         );
  AO22D0 U1400 ( .A1(n206), .A2(n941), .B1(n488), .B2(
        \completionDataOut[7][11] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[11].enDff/theFlop/N3 )
         );
  AO22D0 U1401 ( .A1(n218), .A2(n940), .B1(n925), .B2(
        \completionDataOut[7][23] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[23].enDff/theFlop/N3 )
         );
  AO22D0 U1402 ( .A1(n217), .A2(n940), .B1(n927), .B2(
        \completionDataOut[7][22] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[22].enDff/theFlop/N3 )
         );
  AO22D0 U1403 ( .A1(n219), .A2(n940), .B1(n927), .B2(
        \completionDataOut[7][24] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[24].enDff/theFlop/N3 )
         );
  AO22D0 U1404 ( .A1(n220), .A2(n940), .B1(n925), .B2(
        \completionDataOut[7][25] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[25].enDff/theFlop/N3 )
         );
  AO22D0 U1405 ( .A1(n244), .A2(n933), .B1(n926), .B2(
        \completionDataOut[7][49] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[49].enDff/theFlop/N3 )
         );
  AO22D0 U1406 ( .A1(n201), .A2(n936), .B1(n924), .B2(
        \completionDataOut[7][6] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U1407 ( .A1(n203), .A2(n936), .B1(n924), .B2(
        \completionDataOut[7][8] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U1408 ( .A1(n246), .A2(n933), .B1(n926), .B2(
        \completionDataOut[7][51] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[51].enDff/theFlop/N3 )
         );
  AO22D0 U1409 ( .A1(n204), .A2(n936), .B1(n924), .B2(
        \completionDataOut[7][9] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[9].enDff/theFlop/N3 ) );
  AO22D0 U1410 ( .A1(n243), .A2(n933), .B1(n926), .B2(
        \completionDataOut[7][48] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[48].enDff/theFlop/N3 )
         );
  AO22D0 U1411 ( .A1(n247), .A2(n933), .B1(n926), .B2(
        \completionDataOut[7][52] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[52].enDff/theFlop/N3 )
         );
  AO22D0 U1412 ( .A1(n202), .A2(n936), .B1(n924), .B2(
        \completionDataOut[7][7] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U1413 ( .A1(completionWriteData_i[9]), .A2(n883), .B1(n871), .B2(
        \completionDataOut[5][9] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[9].enDff/theFlop/N3 ) );
  AO22D0 U1414 ( .A1(completionWriteData_i[46]), .A2(n880), .B1(n873), .B2(
        \completionDataOut[5][46] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[46].enDff/theFlop/N3 )
         );
  AO22D0 U1415 ( .A1(completionWriteData_i[43]), .A2(n880), .B1(n873), .B2(
        \completionDataOut[5][43] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[43].enDff/theFlop/N3 )
         );
  AO22D0 U1416 ( .A1(completionWriteData_i[42]), .A2(n880), .B1(n873), .B2(
        \completionDataOut[5][42] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[42].enDff/theFlop/N3 )
         );
  AO22D0 U1417 ( .A1(completionWriteData_i[7]), .A2(n883), .B1(n871), .B2(
        \completionDataOut[5][7] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U1418 ( .A1(completionWriteData_i[8]), .A2(n883), .B1(n871), .B2(
        \completionDataOut[5][8] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U1419 ( .A1(completionWriteData_i[47]), .A2(n880), .B1(n873), .B2(
        \completionDataOut[5][47] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[47].enDff/theFlop/N3 )
         );
  AO22D0 U1420 ( .A1(completionWriteData_i[6]), .A2(n883), .B1(n871), .B2(
        \completionDataOut[5][6] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U1421 ( .A1(n195), .A2(n862), .B1(n836), .B2(
        \completionDataOut[3][0] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U1422 ( .A1(n828), .A2(\completionDataOut[2][5] ), .B1(n809), .B2(
        completionWriteData_i[5]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U1423 ( .A1(n828), .A2(\completionDataOut[2][60] ), .B1(n809), .B2(
        completionWriteData_i[60]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[60].enDff/theFlop/N3 )
         );
  AO22D0 U1424 ( .A1(n834), .A2(\completionDataOut[2][59] ), .B1(n809), .B2(
        completionWriteData_i[59]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[59].enDff/theFlop/N3 )
         );
  AO22D0 U1425 ( .A1(n827), .A2(\completionDataOut[2][69] ), .B1(n808), .B2(
        completionWriteData_i[69]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[69].enDff/theFlop/N3 )
         );
  AO22D0 U1426 ( .A1(n827), .A2(\completionDataOut[2][68] ), .B1(n808), .B2(
        completionWriteData_i[68]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[68].enDff/theFlop/N3 )
         );
  AO22D0 U1427 ( .A1(n828), .A2(\completionDataOut[2][61] ), .B1(n809), .B2(
        completionWriteData_i[61]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[61].enDff/theFlop/N3 )
         );
  AO22D0 U1428 ( .A1(n829), .A2(\completionDataOut[2][51] ), .B1(n810), .B2(
        completionWriteData_i[51]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[51].enDff/theFlop/N3 )
         );
  AO22D0 U1429 ( .A1(n829), .A2(\completionDataOut[2][52] ), .B1(n810), .B2(
        completionWriteData_i[52]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[52].enDff/theFlop/N3 )
         );
  AO22D0 U1430 ( .A1(n215), .A2(n905), .B1(n902), .B2(
        \completionDataOut[6][20] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[20].enDff/theFlop/N3 )
         );
  AO22D0 U1431 ( .A1(n218), .A2(n905), .B1(n899), .B2(
        \completionDataOut[6][23] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[23].enDff/theFlop/N3 )
         );
  AO22D0 U1432 ( .A1(n195), .A2(n904), .B1(n891), .B2(
        \completionDataOut[6][0] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U1433 ( .A1(n209), .A2(n904), .B1(n891), .B2(
        \completionDataOut[6][14] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[14].enDff/theFlop/N3 )
         );
  AO22D0 U1434 ( .A1(n219), .A2(n905), .B1(n901), .B2(
        \completionDataOut[6][24] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[24].enDff/theFlop/N3 )
         );
  AO22D0 U1435 ( .A1(n216), .A2(n905), .B1(n902), .B2(
        \completionDataOut[6][21] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[21].enDff/theFlop/N3 )
         );
  AO22D0 U1436 ( .A1(n205), .A2(n904), .B1(n891), .B2(
        \completionDataOut[6][10] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[10].enDff/theFlop/N3 )
         );
  AO22D0 U1437 ( .A1(n217), .A2(n905), .B1(n901), .B2(
        \completionDataOut[6][22] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[22].enDff/theFlop/N3 )
         );
  AO22D0 U1438 ( .A1(n207), .A2(n904), .B1(n891), .B2(
        \completionDataOut[6][12] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[12].enDff/theFlop/N3 )
         );
  AO22D0 U1439 ( .A1(n206), .A2(n904), .B1(n891), .B2(
        \completionDataOut[6][11] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[11].enDff/theFlop/N3 )
         );
  AO22D0 U1440 ( .A1(n208), .A2(n904), .B1(n891), .B2(
        \completionDataOut[6][13] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[13].enDff/theFlop/N3 )
         );
  AO22D0 U1441 ( .A1(n220), .A2(n905), .B1(n899), .B2(
        \completionDataOut[6][25] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[25].enDff/theFlop/N3 )
         );
  AO22D0 U1442 ( .A1(n224), .A2(n931), .B1(n928), .B2(
        \completionDataOut[7][29] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[29].enDff/theFlop/N3 )
         );
  AO22D0 U1443 ( .A1(n214), .A2(n930), .B1(n917), .B2(
        \completionDataOut[7][19] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[19].enDff/theFlop/N3 )
         );
  AO22D0 U1444 ( .A1(n222), .A2(n931), .B1(n488), .B2(
        \completionDataOut[7][27] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[27].enDff/theFlop/N3 )
         );
  AO22D0 U1445 ( .A1(n210), .A2(n930), .B1(n917), .B2(
        \completionDataOut[7][15] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[15].enDff/theFlop/N3 )
         );
  AO22D0 U1446 ( .A1(n221), .A2(n931), .B1(n488), .B2(
        \completionDataOut[7][26] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[26].enDff/theFlop/N3 )
         );
  AO22D0 U1447 ( .A1(n225), .A2(n931), .B1(n925), .B2(
        \completionDataOut[7][30] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[30].enDff/theFlop/N3 )
         );
  AO22D0 U1448 ( .A1(n197), .A2(n931), .B1(n927), .B2(
        \completionDataOut[7][2] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U1449 ( .A1(n211), .A2(n930), .B1(n917), .B2(
        \completionDataOut[7][16] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[16].enDff/theFlop/N3 )
         );
  AO22D0 U1450 ( .A1(n196), .A2(n930), .B1(n917), .B2(
        \completionDataOut[7][1] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U1451 ( .A1(n212), .A2(n930), .B1(n917), .B2(
        \completionDataOut[7][17] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[17].enDff/theFlop/N3 )
         );
  AO22D0 U1452 ( .A1(n223), .A2(n931), .B1(n928), .B2(
        \completionDataOut[7][28] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[28].enDff/theFlop/N3 )
         );
  AO22D0 U1453 ( .A1(n213), .A2(n930), .B1(n917), .B2(
        \completionDataOut[7][18] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[18].enDff/theFlop/N3 )
         );
  AO22D0 U1454 ( .A1(completionWriteData_i[30]), .A2(n887), .B1(n872), .B2(
        \completionDataOut[5][30] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[30].enDff/theFlop/N3 )
         );
  AO22D0 U1455 ( .A1(completionWriteData_i[2]), .A2(n887), .B1(n874), .B2(
        \completionDataOut[5][2] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U1456 ( .A1(n257), .A2(n911), .B1(n896), .B2(
        \completionDataOut[6][62] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[62].enDff/theFlop/N3 )
         );
  AO22D0 U1457 ( .A1(n256), .A2(n911), .B1(n896), .B2(
        \completionDataOut[6][61] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[61].enDff/theFlop/N3 )
         );
  AO22D0 U1458 ( .A1(n255), .A2(n911), .B1(n896), .B2(
        \completionDataOut[6][60] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[60].enDff/theFlop/N3 )
         );
  AO22D0 U1459 ( .A1(n226), .A2(n906), .B1(n892), .B2(
        \completionDataOut[6][31] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[31].enDff/theFlop/N3 )
         );
  AO22D0 U1460 ( .A1(completionWriteData_i[58]), .A2(n908), .B1(n895), .B2(
        \completionDataOut[6][58] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[58].enDff/theFlop/N3 )
         );
  AO22D0 U1461 ( .A1(n258), .A2(n911), .B1(n896), .B2(
        \completionDataOut[6][63] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[63].enDff/theFlop/N3 )
         );
  AO22D0 U1462 ( .A1(n252), .A2(n908), .B1(n895), .B2(
        \completionDataOut[6][57] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[57].enDff/theFlop/N3 )
         );
  AO22D0 U1463 ( .A1(completionWriteData_i[56]), .A2(n908), .B1(n895), .B2(
        \completionDataOut[6][56] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[56].enDff/theFlop/N3 )
         );
  AO22D0 U1464 ( .A1(n250), .A2(n908), .B1(n895), .B2(
        \completionDataOut[6][55] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[55].enDff/theFlop/N3 )
         );
  AO22D0 U1465 ( .A1(n230), .A2(n906), .B1(n892), .B2(
        \completionDataOut[6][35] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[35].enDff/theFlop/N3 )
         );
  AO22D0 U1466 ( .A1(completionWriteData_i[40]), .A2(n913), .B1(n893), .B2(
        \completionDataOut[6][40] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[40].enDff/theFlop/N3 )
         );
  AO22D0 U1467 ( .A1(n234), .A2(n913), .B1(n893), .B2(
        \completionDataOut[6][39] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[39].enDff/theFlop/N3 )
         );
  AO22D0 U1468 ( .A1(n233), .A2(n913), .B1(n893), .B2(
        \completionDataOut[6][38] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[38].enDff/theFlop/N3 )
         );
  AO22D0 U1469 ( .A1(n232), .A2(n916), .B1(n893), .B2(
        \completionDataOut[6][37] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[37].enDff/theFlop/N3 )
         );
  AO22D0 U1470 ( .A1(n231), .A2(n906), .B1(n892), .B2(
        \completionDataOut[6][36] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[36].enDff/theFlop/N3 )
         );
  AO22D0 U1471 ( .A1(completionWriteData_i[34]), .A2(n906), .B1(n892), .B2(
        \completionDataOut[6][34] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[34].enDff/theFlop/N3 )
         );
  AO22D0 U1472 ( .A1(n249), .A2(n908), .B1(n895), .B2(
        \completionDataOut[6][54] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[54].enDff/theFlop/N3 )
         );
  AO22D0 U1473 ( .A1(completionWriteData_i[33]), .A2(n906), .B1(n892), .B2(
        \completionDataOut[6][33] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[33].enDff/theFlop/N3 )
         );
  AO22D0 U1474 ( .A1(n248), .A2(n908), .B1(n895), .B2(
        \completionDataOut[6][53] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[53].enDff/theFlop/N3 )
         );
  AO22D0 U1475 ( .A1(n198), .A2(n913), .B1(n893), .B2(
        \completionDataOut[6][3] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U1476 ( .A1(n200), .A2(n911), .B1(n896), .B2(
        \completionDataOut[6][5] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U1477 ( .A1(n236), .A2(n913), .B1(n893), .B2(
        \completionDataOut[6][41] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[41].enDff/theFlop/N3 )
         );
  AO22D0 U1478 ( .A1(completionWriteData_i[32]), .A2(n906), .B1(n892), .B2(
        \completionDataOut[6][32] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[32].enDff/theFlop/N3 )
         );
  CKBD1 U1479 ( .I(n1275), .Z(n902) );
  CKBD1 U1480 ( .I(n494), .Z(n916) );
  AO22D0 U1481 ( .A1(completionWriteData_i[12]), .A2(n877), .B1(n871), .B2(
        \completionDataOut[5][12] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[12].enDff/theFlop/N3 )
         );
  AO22D0 U1482 ( .A1(completionWriteData_i[13]), .A2(n877), .B1(n873), .B2(
        \completionDataOut[5][13] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[13].enDff/theFlop/N3 )
         );
  AO22D0 U1483 ( .A1(completionWriteData_i[11]), .A2(n877), .B1(n1271), .B2(
        \completionDataOut[5][11] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[11].enDff/theFlop/N3 )
         );
  AO22D0 U1484 ( .A1(completionWriteData_i[14]), .A2(n877), .B1(n876), .B2(
        \completionDataOut[5][14] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[14].enDff/theFlop/N3 )
         );
  AO22D0 U1485 ( .A1(n216), .A2(n878), .B1(n872), .B2(
        \completionDataOut[5][21] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[21].enDff/theFlop/N3 )
         );
  AO22D0 U1486 ( .A1(completionWriteData_i[24]), .A2(n878), .B1(n874), .B2(
        \completionDataOut[5][24] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[24].enDff/theFlop/N3 )
         );
  AO22D0 U1487 ( .A1(completionWriteData_i[22]), .A2(n878), .B1(n874), .B2(
        \completionDataOut[5][22] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[22].enDff/theFlop/N3 )
         );
  AO22D0 U1488 ( .A1(completionWriteData_i[25]), .A2(n878), .B1(n872), .B2(
        \completionDataOut[5][25] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[25].enDff/theFlop/N3 )
         );
  AO22D0 U1489 ( .A1(completionWriteData_i[0]), .A2(n877), .B1(n1271), .B2(
        \completionDataOut[5][0] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U1490 ( .A1(completionWriteData_i[23]), .A2(n878), .B1(n872), .B2(
        \completionDataOut[5][23] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[23].enDff/theFlop/N3 )
         );
  AO22D0 U1491 ( .A1(n205), .A2(n877), .B1(n1271), .B2(
        \completionDataOut[5][10] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[10].enDff/theFlop/N3 )
         );
  AO22D0 U1492 ( .A1(n215), .A2(n878), .B1(n874), .B2(
        \completionDataOut[5][20] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[20].enDff/theFlop/N3 )
         );
  AO22D0 U1493 ( .A1(n201), .A2(n856), .B1(n843), .B2(
        \completionDataOut[3][6] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U1494 ( .A1(n204), .A2(n856), .B1(n843), .B2(
        \completionDataOut[3][9] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[9].enDff/theFlop/N3 ) );
  AO22D0 U1495 ( .A1(n203), .A2(n856), .B1(n843), .B2(
        \completionDataOut[3][8] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U1496 ( .A1(n202), .A2(n856), .B1(n843), .B2(
        \completionDataOut[3][7] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U1497 ( .A1(n825), .A2(\completionDataOut[2][45] ), .B1(n812), .B2(
        completionWriteData_i[45]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[45].enDff/theFlop/N3 )
         );
  AO22D0 U1498 ( .A1(n826), .A2(\completionDataOut[2][53] ), .B1(n810), .B2(
        completionWriteData_i[53]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[53].enDff/theFlop/N3 )
         );
  AO22D0 U1499 ( .A1(n825), .A2(\completionDataOut[2][42] ), .B1(n812), .B2(
        completionWriteData_i[42]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[42].enDff/theFlop/N3 )
         );
  AO22D0 U1500 ( .A1(n826), .A2(\completionDataOut[2][55] ), .B1(n810), .B2(
        completionWriteData_i[55]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[55].enDff/theFlop/N3 )
         );
  AO22D0 U1501 ( .A1(n826), .A2(\completionDataOut[2][58] ), .B1(n809), .B2(
        completionWriteData_i[58]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[58].enDff/theFlop/N3 )
         );
  AO22D0 U1502 ( .A1(n826), .A2(\completionDataOut[2][54] ), .B1(n810), .B2(
        n249), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[54].enDff/theFlop/N3 )
         );
  AO22D0 U1503 ( .A1(n825), .A2(\completionDataOut[2][44] ), .B1(n812), .B2(
        completionWriteData_i[44]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[44].enDff/theFlop/N3 )
         );
  AO22D0 U1504 ( .A1(n825), .A2(\completionDataOut[2][47] ), .B1(n811), .B2(
        completionWriteData_i[47]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[47].enDff/theFlop/N3 )
         );
  AO22D0 U1505 ( .A1(n826), .A2(\completionDataOut[2][56] ), .B1(n810), .B2(
        completionWriteData_i[56]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[56].enDff/theFlop/N3 )
         );
  AO22D0 U1506 ( .A1(n825), .A2(\completionDataOut[2][46] ), .B1(n811), .B2(
        completionWriteData_i[46]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[46].enDff/theFlop/N3 )
         );
  AO22D0 U1507 ( .A1(n826), .A2(\completionDataOut[2][57] ), .B1(n809), .B2(
        completionWriteData_i[57]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[57].enDff/theFlop/N3 )
         );
  AO22D0 U1508 ( .A1(n825), .A2(\completionDataOut[2][43] ), .B1(n812), .B2(
        completionWriteData_i[43]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[43].enDff/theFlop/N3 )
         );
  AO22D0 U1509 ( .A1(n245), .A2(n853), .B1(n848), .B2(
        \completionDataOut[3][50] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[50].enDff/theFlop/N3 )
         );
  AO22D0 U1510 ( .A1(n244), .A2(n853), .B1(n845), .B2(
        \completionDataOut[3][49] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[49].enDff/theFlop/N3 )
         );
  AO22D0 U1511 ( .A1(n246), .A2(n853), .B1(n845), .B2(
        \completionDataOut[3][51] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[51].enDff/theFlop/N3 )
         );
  AO22D0 U1512 ( .A1(n243), .A2(n853), .B1(n845), .B2(
        \completionDataOut[3][48] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[48].enDff/theFlop/N3 )
         );
  AO22D0 U1513 ( .A1(n247), .A2(n853), .B1(n845), .B2(
        \completionDataOut[3][52] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[52].enDff/theFlop/N3 )
         );
  AO22D0 U1514 ( .A1(n199), .A2(n853), .B1(n848), .B2(
        \completionDataOut[3][4] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U1515 ( .A1(completionWriteData_i[68]), .A2(n909), .B1(n897), .B2(
        \completionDataOut[6][68] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[68].enDff/theFlop/N3 )
         );
  AO22D0 U1516 ( .A1(completionWriteData_i[67]), .A2(n909), .B1(n897), .B2(
        \completionDataOut[6][67] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[67].enDff/theFlop/N3 )
         );
  AO22D0 U1517 ( .A1(completionWriteData_i[66]), .A2(n909), .B1(n897), .B2(
        \completionDataOut[6][66] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[66].enDff/theFlop/N3 )
         );
  AO22D0 U1518 ( .A1(completionWriteData_i[65]), .A2(n909), .B1(n897), .B2(
        \completionDataOut[6][65] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[65].enDff/theFlop/N3 )
         );
  AO22D0 U1519 ( .A1(completionWriteData_i[64]), .A2(n909), .B1(n897), .B2(
        \completionDataOut[6][64] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[64].enDff/theFlop/N3 )
         );
  AO22D0 U1520 ( .A1(n237), .A2(n907), .B1(n894), .B2(
        \completionDataOut[6][42] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[42].enDff/theFlop/N3 )
         );
  AO22D0 U1521 ( .A1(n238), .A2(n907), .B1(n894), .B2(
        \completionDataOut[6][43] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[43].enDff/theFlop/N3 )
         );
  AO22D0 U1522 ( .A1(n239), .A2(n907), .B1(n894), .B2(
        \completionDataOut[6][44] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[44].enDff/theFlop/N3 )
         );
  AO22D0 U1523 ( .A1(n240), .A2(n907), .B1(n894), .B2(
        \completionDataOut[6][45] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[45].enDff/theFlop/N3 )
         );
  AO22D0 U1524 ( .A1(n241), .A2(n907), .B1(n894), .B2(
        \completionDataOut[6][46] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[46].enDff/theFlop/N3 )
         );
  AO22D0 U1525 ( .A1(n242), .A2(n907), .B1(n894), .B2(
        \completionDataOut[6][47] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[47].enDff/theFlop/N3 )
         );
  AO22D0 U1526 ( .A1(completionWriteData_i[69]), .A2(n909), .B1(n897), .B2(
        \completionDataOut[6][69] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[69].enDff/theFlop/N3 )
         );
  CKBD1 U1527 ( .I(n1275), .Z(n903) );
  AO22D0 U1528 ( .A1(n208), .A2(n861), .B1(n836), .B2(
        \completionDataOut[3][13] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[13].enDff/theFlop/N3 )
         );
  AO22D0 U1529 ( .A1(n209), .A2(n861), .B1(n836), .B2(
        \completionDataOut[3][14] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[14].enDff/theFlop/N3 )
         );
  AO22D0 U1530 ( .A1(n207), .A2(n861), .B1(n836), .B2(
        \completionDataOut[3][12] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[12].enDff/theFlop/N3 )
         );
  AO22D0 U1531 ( .A1(n205), .A2(n861), .B1(n836), .B2(
        \completionDataOut[3][10] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[10].enDff/theFlop/N3 )
         );
  AO22D0 U1532 ( .A1(n217), .A2(n860), .B1(n846), .B2(
        \completionDataOut[3][22] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[22].enDff/theFlop/N3 )
         );
  AO22D0 U1533 ( .A1(n220), .A2(n860), .B1(n844), .B2(
        \completionDataOut[3][25] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[25].enDff/theFlop/N3 )
         );
  AO22D0 U1534 ( .A1(n216), .A2(n860), .B1(n847), .B2(
        \completionDataOut[3][21] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[21].enDff/theFlop/N3 )
         );
  AO22D0 U1535 ( .A1(n206), .A2(n861), .B1(n836), .B2(
        \completionDataOut[3][11] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[11].enDff/theFlop/N3 )
         );
  AO22D0 U1536 ( .A1(n218), .A2(n860), .B1(n844), .B2(
        \completionDataOut[3][23] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[23].enDff/theFlop/N3 )
         );
  AO22D0 U1537 ( .A1(n219), .A2(n860), .B1(n846), .B2(
        \completionDataOut[3][24] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[24].enDff/theFlop/N3 )
         );
  AO22D0 U1538 ( .A1(n830), .A2(\completionDataOut[2][38] ), .B1(n818), .B2(
        completionWriteData_i[38]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[38].enDff/theFlop/N3 )
         );
  AO22D0 U1539 ( .A1(n823), .A2(\completionDataOut[2][24] ), .B1(n817), .B2(
        completionWriteData_i[24]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[24].enDff/theFlop/N3 )
         );
  AO22D0 U1540 ( .A1(n823), .A2(\completionDataOut[2][25] ), .B1(n817), .B2(
        completionWriteData_i[25]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[25].enDff/theFlop/N3 )
         );
  AO22D0 U1541 ( .A1(n830), .A2(\completionDataOut[2][39] ), .B1(n818), .B2(
        completionWriteData_i[39]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[39].enDff/theFlop/N3 )
         );
  AO22D0 U1542 ( .A1(n831), .A2(\completionDataOut[2][27] ), .B1(n817), .B2(
        completionWriteData_i[27]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[27].enDff/theFlop/N3 )
         );
  AO22D0 U1543 ( .A1(n831), .A2(\completionDataOut[2][28] ), .B1(n817), .B2(
        completionWriteData_i[28]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[28].enDff/theFlop/N3 )
         );
  AO22D0 U1544 ( .A1(n824), .A2(\completionDataOut[2][35] ), .B1(n818), .B2(
        completionWriteData_i[35]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[35].enDff/theFlop/N3 )
         );
  AO22D0 U1545 ( .A1(n824), .A2(\completionDataOut[2][36] ), .B1(n818), .B2(
        completionWriteData_i[36]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[36].enDff/theFlop/N3 )
         );
  AO22D0 U1546 ( .A1(n833), .A2(\completionDataOut[2][26] ), .B1(n817), .B2(
        completionWriteData_i[26]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[26].enDff/theFlop/N3 )
         );
  AO22D0 U1547 ( .A1(n833), .A2(\completionDataOut[2][37] ), .B1(n818), .B2(
        completionWriteData_i[37]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[37].enDff/theFlop/N3 )
         );
  AO22D0 U1548 ( .A1(n229), .A2(n939), .B1(n918), .B2(
        \completionDataOut[7][34] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[34].enDff/theFlop/N3 )
         );
  AO22D0 U1549 ( .A1(n250), .A2(n937), .B1(n921), .B2(
        \completionDataOut[7][55] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[55].enDff/theFlop/N3 )
         );
  AO22D0 U1550 ( .A1(n251), .A2(n937), .B1(n921), .B2(
        \completionDataOut[7][56] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[56].enDff/theFlop/N3 )
         );
  AO22D0 U1551 ( .A1(n252), .A2(n937), .B1(n921), .B2(
        \completionDataOut[7][57] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[57].enDff/theFlop/N3 )
         );
  AO22D0 U1552 ( .A1(n234), .A2(n932), .B1(n919), .B2(
        \completionDataOut[7][39] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[39].enDff/theFlop/N3 )
         );
  AO22D0 U1553 ( .A1(n198), .A2(n932), .B1(n919), .B2(
        \completionDataOut[7][3] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U1554 ( .A1(n200), .A2(n934), .B1(n922), .B2(
        \completionDataOut[7][5] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U1555 ( .A1(n254), .A2(n934), .B1(n922), .B2(
        \completionDataOut[7][59] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[59].enDff/theFlop/N3 )
         );
  AO22D0 U1556 ( .A1(n253), .A2(n937), .B1(n921), .B2(
        \completionDataOut[7][58] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[58].enDff/theFlop/N3 )
         );
  AO22D0 U1557 ( .A1(n226), .A2(n942), .B1(n918), .B2(
        \completionDataOut[7][31] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[31].enDff/theFlop/N3 )
         );
  AO22D0 U1558 ( .A1(n227), .A2(n939), .B1(n918), .B2(
        \completionDataOut[7][32] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[32].enDff/theFlop/N3 )
         );
  AO22D0 U1559 ( .A1(n228), .A2(n939), .B1(n918), .B2(
        \completionDataOut[7][33] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[33].enDff/theFlop/N3 )
         );
  AO22D0 U1560 ( .A1(n255), .A2(n934), .B1(n922), .B2(
        \completionDataOut[7][60] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[60].enDff/theFlop/N3 )
         );
  AO22D0 U1561 ( .A1(n230), .A2(n939), .B1(n918), .B2(
        \completionDataOut[7][35] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[35].enDff/theFlop/N3 )
         );
  AO22D0 U1562 ( .A1(n231), .A2(n939), .B1(n918), .B2(
        \completionDataOut[7][36] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[36].enDff/theFlop/N3 )
         );
  AO22D0 U1563 ( .A1(n232), .A2(n932), .B1(n919), .B2(
        \completionDataOut[7][37] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[37].enDff/theFlop/N3 )
         );
  AO22D0 U1564 ( .A1(n233), .A2(n932), .B1(n919), .B2(
        \completionDataOut[7][38] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[38].enDff/theFlop/N3 )
         );
  AO22D0 U1565 ( .A1(n256), .A2(n934), .B1(n922), .B2(
        \completionDataOut[7][61] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[61].enDff/theFlop/N3 )
         );
  AO22D0 U1566 ( .A1(n235), .A2(n932), .B1(n919), .B2(
        \completionDataOut[7][40] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[40].enDff/theFlop/N3 )
         );
  AO22D0 U1567 ( .A1(completionWriteData_i[54]), .A2(n937), .B1(n921), .B2(
        \completionDataOut[7][54] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[54].enDff/theFlop/N3 )
         );
  AO22D0 U1568 ( .A1(n236), .A2(n932), .B1(n919), .B2(
        \completionDataOut[7][41] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[41].enDff/theFlop/N3 )
         );
  CKBD1 U1569 ( .I(n943), .Z(n942) );
  AO22D0 U1570 ( .A1(n258), .A2(n934), .B1(n922), .B2(
        \completionDataOut[7][63] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[63].enDff/theFlop/N3 )
         );
  AO22D0 U1571 ( .A1(n257), .A2(n934), .B1(n922), .B2(
        \completionDataOut[7][62] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[62].enDff/theFlop/N3 )
         );
  CKBD1 U1572 ( .I(n488), .Z(n928) );
  AO22D0 U1573 ( .A1(completionWriteData_i[4]), .A2(n885), .B1(n867), .B2(
        \completionDataOut[5][4] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U1574 ( .A1(completionWriteData_i[49]), .A2(n885), .B1(n867), .B2(
        \completionDataOut[5][49] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[49].enDff/theFlop/N3 )
         );
  AO22D0 U1575 ( .A1(n262), .A2(n882), .B1(n870), .B2(
        \completionDataOut[5][67] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[67].enDff/theFlop/N3 )
         );
  AO22D0 U1576 ( .A1(n264), .A2(n882), .B1(n870), .B2(
        \completionDataOut[5][69] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[69].enDff/theFlop/N3 )
         );
  AO22D0 U1577 ( .A1(n259), .A2(n882), .B1(n870), .B2(
        \completionDataOut[5][64] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[64].enDff/theFlop/N3 )
         );
  AO22D0 U1578 ( .A1(n263), .A2(n882), .B1(n870), .B2(
        \completionDataOut[5][68] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[68].enDff/theFlop/N3 )
         );
  AO22D0 U1579 ( .A1(n261), .A2(n882), .B1(n870), .B2(
        \completionDataOut[5][66] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[66].enDff/theFlop/N3 )
         );
  AO22D0 U1580 ( .A1(completionWriteData_i[50]), .A2(n885), .B1(n867), .B2(
        \completionDataOut[5][50] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[50].enDff/theFlop/N3 )
         );
  AO22D0 U1581 ( .A1(completionWriteData_i[52]), .A2(n885), .B1(n867), .B2(
        \completionDataOut[5][52] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[52].enDff/theFlop/N3 )
         );
  AO22D0 U1582 ( .A1(n260), .A2(n882), .B1(n870), .B2(
        \completionDataOut[5][65] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[65].enDff/theFlop/N3 )
         );
  AO22D0 U1583 ( .A1(completionWriteData_i[51]), .A2(n885), .B1(n867), .B2(
        \completionDataOut[5][51] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[51].enDff/theFlop/N3 )
         );
  CKBD1 U1584 ( .I(n1271), .Z(n876) );
  AO22D0 U1585 ( .A1(n239), .A2(n938), .B1(n920), .B2(
        \completionDataOut[7][44] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[44].enDff/theFlop/N3 )
         );
  AO22D0 U1586 ( .A1(n240), .A2(n938), .B1(n920), .B2(
        \completionDataOut[7][45] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[45].enDff/theFlop/N3 )
         );
  AO22D0 U1587 ( .A1(n241), .A2(n938), .B1(n920), .B2(
        \completionDataOut[7][46] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[46].enDff/theFlop/N3 )
         );
  AO22D0 U1588 ( .A1(n238), .A2(n938), .B1(n920), .B2(
        \completionDataOut[7][43] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[43].enDff/theFlop/N3 )
         );
  AO22D0 U1589 ( .A1(n260), .A2(n935), .B1(n923), .B2(
        \completionDataOut[7][65] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[65].enDff/theFlop/N3 )
         );
  AO22D0 U1590 ( .A1(n259), .A2(n935), .B1(n923), .B2(
        \completionDataOut[7][64] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[64].enDff/theFlop/N3 )
         );
  AO22D0 U1591 ( .A1(n261), .A2(n935), .B1(n923), .B2(
        \completionDataOut[7][66] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[66].enDff/theFlop/N3 )
         );
  AO22D0 U1592 ( .A1(n262), .A2(n935), .B1(n923), .B2(
        \completionDataOut[7][67] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[67].enDff/theFlop/N3 )
         );
  AO22D0 U1593 ( .A1(n264), .A2(n935), .B1(n923), .B2(
        \completionDataOut[7][69] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[69].enDff/theFlop/N3 )
         );
  AO22D0 U1594 ( .A1(n263), .A2(n935), .B1(n923), .B2(
        \completionDataOut[7][68] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[68].enDff/theFlop/N3 )
         );
  AO22D0 U1595 ( .A1(n242), .A2(n938), .B1(n920), .B2(
        \completionDataOut[7][47] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[47].enDff/theFlop/N3 )
         );
  CKBD1 U1596 ( .I(n488), .Z(n929) );
  CKBD1 U1597 ( .I(n1280), .Z(n943) );
  AO22D0 U1598 ( .A1(completionWriteData_i[55]), .A2(n881), .B1(n868), .B2(
        \completionDataOut[5][55] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[55].enDff/theFlop/N3 )
         );
  AO22D0 U1599 ( .A1(completionWriteData_i[53]), .A2(n881), .B1(n868), .B2(
        \completionDataOut[5][53] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[53].enDff/theFlop/N3 )
         );
  AO22D0 U1600 ( .A1(completionWriteData_i[54]), .A2(n881), .B1(n868), .B2(
        \completionDataOut[5][54] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[54].enDff/theFlop/N3 )
         );
  AO22D0 U1601 ( .A1(n251), .A2(n881), .B1(n868), .B2(
        \completionDataOut[5][56] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[56].enDff/theFlop/N3 )
         );
  AO22D0 U1602 ( .A1(n258), .A2(n884), .B1(n869), .B2(
        \completionDataOut[5][63] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[63].enDff/theFlop/N3 )
         );
  AO22D0 U1603 ( .A1(completionWriteData_i[62]), .A2(n884), .B1(n869), .B2(
        \completionDataOut[5][62] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[62].enDff/theFlop/N3 )
         );
  AO22D0 U1604 ( .A1(completionWriteData_i[61]), .A2(n884), .B1(n869), .B2(
        \completionDataOut[5][61] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[61].enDff/theFlop/N3 )
         );
  AO22D0 U1605 ( .A1(completionWriteData_i[60]), .A2(n884), .B1(n869), .B2(
        \completionDataOut[5][60] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[60].enDff/theFlop/N3 )
         );
  AO22D0 U1606 ( .A1(n253), .A2(n881), .B1(n868), .B2(
        \completionDataOut[5][58] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[58].enDff/theFlop/N3 )
         );
  AO22D0 U1607 ( .A1(n252), .A2(n881), .B1(n868), .B2(
        \completionDataOut[5][57] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[57].enDff/theFlop/N3 )
         );
  AO22D0 U1608 ( .A1(n228), .A2(n879), .B1(n865), .B2(
        \completionDataOut[5][33] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[33].enDff/theFlop/N3 )
         );
  AO22D0 U1609 ( .A1(completionWriteData_i[39]), .A2(n886), .B1(n866), .B2(
        \completionDataOut[5][39] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[39].enDff/theFlop/N3 )
         );
  AO22D0 U1610 ( .A1(n227), .A2(n879), .B1(n865), .B2(
        \completionDataOut[5][32] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[32].enDff/theFlop/N3 )
         );
  AO22D0 U1611 ( .A1(completionWriteData_i[41]), .A2(n886), .B1(n866), .B2(
        \completionDataOut[5][41] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[41].enDff/theFlop/N3 )
         );
  AO22D0 U1612 ( .A1(n235), .A2(n886), .B1(n866), .B2(
        \completionDataOut[5][40] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[40].enDff/theFlop/N3 )
         );
  AO22D0 U1613 ( .A1(completionWriteData_i[35]), .A2(n879), .B1(n865), .B2(
        \completionDataOut[5][35] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[35].enDff/theFlop/N3 )
         );
  AO22D0 U1614 ( .A1(completionWriteData_i[38]), .A2(n886), .B1(n866), .B2(
        \completionDataOut[5][38] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[38].enDff/theFlop/N3 )
         );
  AO22D0 U1615 ( .A1(completionWriteData_i[37]), .A2(n889), .B1(n866), .B2(
        \completionDataOut[5][37] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[37].enDff/theFlop/N3 )
         );
  AO22D0 U1616 ( .A1(completionWriteData_i[36]), .A2(n879), .B1(n865), .B2(
        \completionDataOut[5][36] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[36].enDff/theFlop/N3 )
         );
  AO22D0 U1617 ( .A1(completionWriteData_i[31]), .A2(n879), .B1(n865), .B2(
        \completionDataOut[5][31] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[31].enDff/theFlop/N3 )
         );
  AO22D0 U1618 ( .A1(n229), .A2(n879), .B1(n865), .B2(
        \completionDataOut[5][34] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[34].enDff/theFlop/N3 )
         );
  AO22D0 U1619 ( .A1(completionWriteData_i[5]), .A2(n884), .B1(n869), .B2(
        \completionDataOut[5][5] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U1620 ( .A1(completionWriteData_i[3]), .A2(n886), .B1(n866), .B2(
        \completionDataOut[5][3] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[3].enDff/theFlop/N3 ) );
  CKBD1 U1621 ( .I(n1271), .Z(n875) );
  CKBD1 U1622 ( .I(n890), .Z(n889) );
  CKBD1 U1623 ( .I(n1272), .Z(n890) );
  NR2D1 U1624 ( .A1(completionWriteAddr_i[1]), .A2(n1269), .ZN(n1303) );
  INVD1 U1625 ( .I(n1304), .ZN(n1278) );
  AO22D0 U1626 ( .A1(n257), .A2(n854), .B1(n841), .B2(
        \completionDataOut[3][62] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[62].enDff/theFlop/N3 )
         );
  AO22D0 U1627 ( .A1(n250), .A2(n857), .B1(n840), .B2(
        \completionDataOut[3][55] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[55].enDff/theFlop/N3 )
         );
  AO22D0 U1628 ( .A1(n255), .A2(n854), .B1(n841), .B2(
        \completionDataOut[3][60] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[60].enDff/theFlop/N3 )
         );
  AO22D0 U1629 ( .A1(n249), .A2(n857), .B1(n840), .B2(
        \completionDataOut[3][54] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[54].enDff/theFlop/N3 )
         );
  AO22D0 U1630 ( .A1(n253), .A2(n857), .B1(n840), .B2(
        \completionDataOut[3][58] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[58].enDff/theFlop/N3 )
         );
  AO22D0 U1631 ( .A1(n254), .A2(n854), .B1(n841), .B2(
        \completionDataOut[3][59] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[59].enDff/theFlop/N3 )
         );
  AO22D0 U1632 ( .A1(n227), .A2(n859), .B1(n837), .B2(
        \completionDataOut[3][32] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[32].enDff/theFlop/N3 )
         );
  AO22D0 U1633 ( .A1(completionWriteData_i[57]), .A2(n857), .B1(n840), .B2(
        \completionDataOut[3][57] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[57].enDff/theFlop/N3 )
         );
  AO22D0 U1634 ( .A1(n229), .A2(n859), .B1(n837), .B2(
        \completionDataOut[3][34] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[34].enDff/theFlop/N3 )
         );
  AO22D0 U1635 ( .A1(completionWriteData_i[63]), .A2(n854), .B1(n841), .B2(
        \completionDataOut[3][63] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[63].enDff/theFlop/N3 )
         );
  AO22D0 U1636 ( .A1(n200), .A2(n854), .B1(n841), .B2(
        \completionDataOut[3][5] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U1637 ( .A1(n226), .A2(n862), .B1(n837), .B2(
        \completionDataOut[3][31] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[31].enDff/theFlop/N3 )
         );
  AO22D0 U1638 ( .A1(n251), .A2(n857), .B1(n840), .B2(
        \completionDataOut[3][56] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[56].enDff/theFlop/N3 )
         );
  AO22D0 U1639 ( .A1(n228), .A2(n859), .B1(n837), .B2(
        \completionDataOut[3][33] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[33].enDff/theFlop/N3 )
         );
  AO22D0 U1640 ( .A1(n231), .A2(n859), .B1(n837), .B2(
        \completionDataOut[3][36] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[36].enDff/theFlop/N3 )
         );
  AO22D0 U1641 ( .A1(n256), .A2(n854), .B1(n841), .B2(
        \completionDataOut[3][61] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[61].enDff/theFlop/N3 )
         );
  AO22D0 U1642 ( .A1(n230), .A2(n859), .B1(n837), .B2(
        \completionDataOut[3][35] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[35].enDff/theFlop/N3 )
         );
  AO22D0 U1643 ( .A1(n240), .A2(n858), .B1(n839), .B2(
        \completionDataOut[3][45] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[45].enDff/theFlop/N3 )
         );
  AO22D0 U1644 ( .A1(n260), .A2(n855), .B1(n842), .B2(
        \completionDataOut[3][65] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[65].enDff/theFlop/N3 )
         );
  AO22D0 U1645 ( .A1(n238), .A2(n858), .B1(n839), .B2(
        \completionDataOut[3][43] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[43].enDff/theFlop/N3 )
         );
  AO22D0 U1646 ( .A1(n263), .A2(n855), .B1(n842), .B2(
        \completionDataOut[3][68] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[68].enDff/theFlop/N3 )
         );
  AO22D0 U1647 ( .A1(n262), .A2(n855), .B1(n842), .B2(
        \completionDataOut[3][67] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[67].enDff/theFlop/N3 )
         );
  AO22D0 U1648 ( .A1(n241), .A2(n858), .B1(n839), .B2(
        \completionDataOut[3][46] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[46].enDff/theFlop/N3 )
         );
  AO22D0 U1649 ( .A1(n261), .A2(n855), .B1(n842), .B2(
        \completionDataOut[3][66] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[66].enDff/theFlop/N3 )
         );
  AO22D0 U1650 ( .A1(n242), .A2(n858), .B1(n839), .B2(
        \completionDataOut[3][47] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[47].enDff/theFlop/N3 )
         );
  AO22D0 U1651 ( .A1(n264), .A2(n855), .B1(n842), .B2(
        \completionDataOut[3][69] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[69].enDff/theFlop/N3 )
         );
  AO22D0 U1652 ( .A1(n239), .A2(n858), .B1(n839), .B2(
        \completionDataOut[3][44] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[44].enDff/theFlop/N3 )
         );
  AO22D0 U1653 ( .A1(n259), .A2(n855), .B1(n842), .B2(
        \completionDataOut[3][64] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[64].enDff/theFlop/N3 )
         );
  AO22D0 U1654 ( .A1(n233), .A2(n852), .B1(n838), .B2(
        \completionDataOut[3][38] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[38].enDff/theFlop/N3 )
         );
  AO22D0 U1655 ( .A1(n234), .A2(n852), .B1(n838), .B2(
        \completionDataOut[3][39] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[39].enDff/theFlop/N3 )
         );
  AO22D0 U1656 ( .A1(n198), .A2(n852), .B1(n838), .B2(
        \completionDataOut[3][3] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U1657 ( .A1(n232), .A2(n852), .B1(n838), .B2(
        \completionDataOut[3][37] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[37].enDff/theFlop/N3 )
         );
  AO22D0 U1658 ( .A1(n196), .A2(n850), .B1(n845), .B2(
        \completionDataOut[3][1] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U1659 ( .A1(n235), .A2(n852), .B1(n838), .B2(
        \completionDataOut[3][40] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[40].enDff/theFlop/N3 )
         );
  AO22D0 U1660 ( .A1(n210), .A2(n850), .B1(n843), .B2(
        \completionDataOut[3][15] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[15].enDff/theFlop/N3 )
         );
  AO22D0 U1661 ( .A1(n236), .A2(n852), .B1(n838), .B2(
        \completionDataOut[3][41] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[41].enDff/theFlop/N3 )
         );
  AO22D0 U1662 ( .A1(n212), .A2(n850), .B1(n848), .B2(
        \completionDataOut[3][17] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[17].enDff/theFlop/N3 )
         );
  AO22D0 U1663 ( .A1(n213), .A2(n850), .B1(n849), .B2(
        \completionDataOut[3][18] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[18].enDff/theFlop/N3 )
         );
  AO22D0 U1664 ( .A1(n214), .A2(n850), .B1(n844), .B2(
        \completionDataOut[3][19] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[19].enDff/theFlop/N3 )
         );
  AO22D0 U1665 ( .A1(n211), .A2(n850), .B1(n849), .B2(
        \completionDataOut[3][16] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[16].enDff/theFlop/N3 )
         );
  CKBD1 U1666 ( .I(n849), .Z(n848) );
  AO22D0 U1667 ( .A1(n197), .A2(n851), .B1(n846), .B2(
        \completionDataOut[3][2] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U1668 ( .A1(n221), .A2(n851), .B1(n849), .B2(
        \completionDataOut[3][26] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[26].enDff/theFlop/N3 )
         );
  AO22D0 U1669 ( .A1(n222), .A2(n851), .B1(n849), .B2(
        \completionDataOut[3][27] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[27].enDff/theFlop/N3 )
         );
  AO22D0 U1670 ( .A1(n223), .A2(n851), .B1(n847), .B2(
        \completionDataOut[3][28] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[28].enDff/theFlop/N3 )
         );
  AO22D0 U1671 ( .A1(n224), .A2(n851), .B1(n847), .B2(
        \completionDataOut[3][29] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[29].enDff/theFlop/N3 )
         );
  AO22D0 U1672 ( .A1(n225), .A2(n851), .B1(n844), .B2(
        \completionDataOut[3][30] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[30].enDff/theFlop/N3 )
         );
  CKBD1 U1673 ( .I(n849), .Z(n847) );
  CKBD1 U1674 ( .I(n1267), .Z(n849) );
  CKBD1 U1675 ( .I(n863), .Z(n862) );
  CKBD1 U1676 ( .I(n1268), .Z(n863) );
  AO22D0 U1677 ( .A1(n822), .A2(\completionDataOut[2][0] ), .B1(
        completionWriteData_i[0]), .B2(n816), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U1678 ( .A1(n827), .A2(\completionDataOut[2][65] ), .B1(n816), .B2(
        completionWriteData_i[65]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[65].enDff/theFlop/N3 )
         );
  AO22D0 U1679 ( .A1(n822), .A2(\completionDataOut[2][10] ), .B1(n816), .B2(
        completionWriteData_i[10]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[10].enDff/theFlop/N3 )
         );
  AO22D0 U1680 ( .A1(n822), .A2(\completionDataOut[2][11] ), .B1(n816), .B2(
        completionWriteData_i[11]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[11].enDff/theFlop/N3 )
         );
  AO22D0 U1681 ( .A1(n822), .A2(\completionDataOut[2][12] ), .B1(n816), .B2(
        completionWriteData_i[12]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[12].enDff/theFlop/N3 )
         );
  AO22D0 U1682 ( .A1(n823), .A2(\completionDataOut[2][21] ), .B1(n814), .B2(
        completionWriteData_i[21]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[21].enDff/theFlop/N3 )
         );
  AO22D0 U1683 ( .A1(n824), .A2(\completionDataOut[2][31] ), .B1(n813), .B2(
        completionWriteData_i[31]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[31].enDff/theFlop/N3 )
         );
  AO22D0 U1684 ( .A1(n823), .A2(\completionDataOut[2][22] ), .B1(n814), .B2(
        completionWriteData_i[22]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[22].enDff/theFlop/N3 )
         );
  AO22D0 U1685 ( .A1(n832), .A2(\completionDataOut[2][1] ), .B1(n814), .B2(
        completionWriteData_i[1]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U1686 ( .A1(n824), .A2(\completionDataOut[2][34] ), .B1(n813), .B2(
        completionWriteData_i[34]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[34].enDff/theFlop/N3 )
         );
  AO22D0 U1687 ( .A1(n832), .A2(\completionDataOut[2][19] ), .B1(n814), .B2(
        completionWriteData_i[19]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[19].enDff/theFlop/N3 )
         );
  AO22D0 U1688 ( .A1(n823), .A2(\completionDataOut[2][20] ), .B1(n814), .B2(
        completionWriteData_i[20]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[20].enDff/theFlop/N3 )
         );
  AO22D0 U1689 ( .A1(n831), .A2(\completionDataOut[2][2] ), .B1(n813), .B2(
        completionWriteData_i[2]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U1690 ( .A1(n831), .A2(\completionDataOut[2][30] ), .B1(n813), .B2(
        completionWriteData_i[30]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[30].enDff/theFlop/N3 )
         );
  AO22D0 U1691 ( .A1(n824), .A2(\completionDataOut[2][32] ), .B1(n813), .B2(
        completionWriteData_i[32]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[32].enDff/theFlop/N3 )
         );
  AO22D0 U1692 ( .A1(n823), .A2(\completionDataOut[2][23] ), .B1(n814), .B2(
        completionWriteData_i[23]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[23].enDff/theFlop/N3 )
         );
  AO22D0 U1693 ( .A1(n824), .A2(\completionDataOut[2][33] ), .B1(n813), .B2(
        completionWriteData_i[33]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[33].enDff/theFlop/N3 )
         );
  AO22D0 U1694 ( .A1(n822), .A2(\completionDataOut[2][13] ), .B1(n815), .B2(
        completionWriteData_i[13]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[13].enDff/theFlop/N3 )
         );
  AO22D0 U1695 ( .A1(n822), .A2(\completionDataOut[2][14] ), .B1(n815), .B2(
        completionWriteData_i[14]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[14].enDff/theFlop/N3 )
         );
  AO22D0 U1696 ( .A1(n832), .A2(\completionDataOut[2][18] ), .B1(n815), .B2(
        completionWriteData_i[18]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[18].enDff/theFlop/N3 )
         );
  AO22D0 U1697 ( .A1(n832), .A2(\completionDataOut[2][16] ), .B1(n815), .B2(
        completionWriteData_i[16]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[16].enDff/theFlop/N3 )
         );
  AO22D0 U1698 ( .A1(n832), .A2(\completionDataOut[2][17] ), .B1(n815), .B2(
        completionWriteData_i[17]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[17].enDff/theFlop/N3 )
         );
  AO22D0 U1699 ( .A1(n833), .A2(\completionDataOut[2][15] ), .B1(n815), .B2(
        completionWriteData_i[15]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[15].enDff/theFlop/N3 )
         );
  CKBD1 U1700 ( .I(n821), .Z(n820) );
  CKBD1 U1701 ( .I(n1264), .Z(n821) );
  CKBD1 U1702 ( .I(n835), .Z(n833) );
  CKBD1 U1703 ( .I(n1265), .Z(n835) );
  NR2D1 U1704 ( .A1(n1302), .A2(n1273), .ZN(n1263) );
  ND2D1 U1705 ( .A1(completionWriteAddr_i[1]), .A2(n1269), .ZN(n1273) );
  IND2D1 U1706 ( .A1(completionWriteAddr_i[2]), .B1(completionWriteEn_i), .ZN(
        n1302) );
  INR2D1 U1707 ( .A1(n1300), .B1(n1299), .ZN(n6) );
  AO22D0 U1708 ( .A1(decodeWriteData_i[4]), .A2(n313), .B1(n504), .B2(
        \managementDataOut[7][4] ), .Z(
        \eachManagementReg[7].managementReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U1709 ( .A1(decodeWriteData_i[5]), .A2(n313), .B1(n504), .B2(
        \managementDataOut[7][5] ), .Z(
        \eachManagementReg[7].managementReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U1710 ( .A1(decodeWriteData_i[1]), .A2(n314), .B1(n504), .B2(
        \managementDataOut[7][1] ), .Z(
        \eachManagementReg[7].managementReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U1711 ( .A1(decodeWriteData_i[8]), .A2(n314), .B1(n504), .B2(
        \managementDataOut[7][8] ), .Z(
        \eachManagementReg[7].managementReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U1712 ( .A1(decodeWriteData_i[6]), .A2(n314), .B1(n504), .B2(
        \managementDataOut[7][6] ), .Z(
        \eachManagementReg[7].managementReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U1713 ( .A1(decodeWriteData_i[3]), .A2(n314), .B1(n505), .B2(
        \managementDataOut[7][3] ), .Z(
        \eachManagementReg[7].managementReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U1714 ( .A1(n272), .A2(n313), .B1(n505), .B2(
        \managementDataOut[7][7] ), .Z(
        \eachManagementReg[7].managementReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U1715 ( .A1(decodeWriteData_i[2]), .A2(n313), .B1(n505), .B2(
        \managementDataOut[7][2] ), .Z(
        \eachManagementReg[7].managementReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U1716 ( .A1(n265), .A2(n313), .B1(n505), .B2(
        \managementDataOut[7][0] ), .Z(
        \eachManagementReg[7].managementReg/eachEnDff[0].enDff/theFlop/N3 ) );
  ND3D1 U1717 ( .A1(decodeWriteAddr_i[0]), .A2(n194), .A3(n1296), .ZN(n1295)
         );
  AO22D0 U1718 ( .A1(n271), .A2(n317), .B1(n502), .B2(
        \managementDataOut[3][6] ), .Z(
        \eachManagementReg[3].managementReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U1719 ( .A1(n270), .A2(n317), .B1(n502), .B2(
        \managementDataOut[3][5] ), .Z(
        \eachManagementReg[3].managementReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U1720 ( .A1(n273), .A2(n318), .B1(n502), .B2(
        \managementDataOut[3][8] ), .Z(
        \eachManagementReg[3].managementReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U1721 ( .A1(decodeWriteData_i[0]), .A2(n318), .B1(n502), .B2(
        \managementDataOut[3][0] ), .Z(
        \eachManagementReg[3].managementReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U1722 ( .A1(n269), .A2(n318), .B1(n502), .B2(
        \managementDataOut[3][4] ), .Z(
        \eachManagementReg[3].managementReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U1723 ( .A1(n267), .A2(n318), .B1(n503), .B2(
        \managementDataOut[3][2] ), .Z(
        \eachManagementReg[3].managementReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U1724 ( .A1(n268), .A2(n317), .B1(n503), .B2(
        \managementDataOut[3][3] ), .Z(
        \eachManagementReg[3].managementReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U1725 ( .A1(n266), .A2(n317), .B1(n503), .B2(
        \managementDataOut[3][1] ), .Z(
        \eachManagementReg[3].managementReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U1726 ( .A1(n272), .A2(n317), .B1(n503), .B2(
        \managementDataOut[3][7] ), .Z(
        \eachManagementReg[3].managementReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U1727 ( .A1(n267), .A2(n316), .B1(n807), .B2(
        \managementDataOut[5][2] ), .Z(
        \eachManagementReg[5].managementReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U1728 ( .A1(n270), .A2(n315), .B1(n807), .B2(
        \managementDataOut[5][5] ), .Z(
        \eachManagementReg[5].managementReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U1729 ( .A1(n271), .A2(n315), .B1(n807), .B2(
        \managementDataOut[5][6] ), .Z(
        \eachManagementReg[5].managementReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U1730 ( .A1(n268), .A2(n316), .B1(n807), .B2(
        \managementDataOut[5][3] ), .Z(
        \eachManagementReg[5].managementReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U1731 ( .A1(n269), .A2(n316), .B1(n807), .B2(
        \managementDataOut[5][4] ), .Z(
        \eachManagementReg[5].managementReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U1732 ( .A1(n273), .A2(n316), .B1(n1289), .B2(
        \managementDataOut[5][8] ), .Z(
        \eachManagementReg[5].managementReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U1733 ( .A1(n265), .A2(n315), .B1(n1289), .B2(
        \managementDataOut[5][0] ), .Z(
        \eachManagementReg[5].managementReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U1734 ( .A1(decodeWriteData_i[7]), .A2(n315), .B1(n1289), .B2(
        \managementDataOut[5][7] ), .Z(
        \eachManagementReg[5].managementReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U1735 ( .A1(n266), .A2(n315), .B1(n1289), .B2(
        \managementDataOut[5][1] ), .Z(
        \eachManagementReg[5].managementReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AOI22D1 U1736 ( .A1(n1082), .A2(\completionDataOut[1][63] ), .B1(n1083), 
        .B2(\completionDataOut[3][63] ), .ZN(n1815) );
  AOI22D1 U1737 ( .A1(n492), .A2(\completionDataOut[0][63] ), .B1(n1057), .B2(
        \completionDataOut[2][63] ), .ZN(n1814) );
  AOI22D1 U1738 ( .A1(n1227), .A2(\completionDataOut[5][18] ), .B1(n1239), 
        .B2(\completionDataOut[7][18] ), .ZN(n1897) );
  AOI22D1 U1739 ( .A1(n1202), .A2(\completionDataOut[4][18] ), .B1(n1214), 
        .B2(\completionDataOut[6][18] ), .ZN(n1896) );
  AOI22D1 U1740 ( .A1(n1176), .A2(\completionDataOut[1][18] ), .B1(n1189), 
        .B2(\completionDataOut[3][18] ), .ZN(n1895) );
  AOI22D1 U1741 ( .A1(n1151), .A2(\completionDataOut[0][18] ), .B1(n1163), 
        .B2(\completionDataOut[2][18] ), .ZN(n1894) );
  AOI22D1 U1742 ( .A1(n1176), .A2(\completionDataOut[1][17] ), .B1(n1189), 
        .B2(\completionDataOut[3][17] ), .ZN(n1893) );
  AOI22D1 U1743 ( .A1(n1151), .A2(\completionDataOut[0][17] ), .B1(n1163), 
        .B2(\completionDataOut[2][17] ), .ZN(n1892) );
  AOI22D1 U1744 ( .A1(n1179), .A2(\completionDataOut[1][16] ), .B1(n1196), 
        .B2(\completionDataOut[3][16] ), .ZN(n1889) );
  AOI22D1 U1745 ( .A1(n1154), .A2(\completionDataOut[0][16] ), .B1(n1170), 
        .B2(\completionDataOut[2][16] ), .ZN(n1888) );
  AOI22D1 U1746 ( .A1(n1082), .A2(\completionDataOut[1][64] ), .B1(n1083), 
        .B2(\completionDataOut[3][64] ), .ZN(n1819) );
  AOI22D1 U1747 ( .A1(n492), .A2(\completionDataOut[0][64] ), .B1(n1057), .B2(
        \completionDataOut[2][64] ), .ZN(n1818) );
  AOI22D1 U1748 ( .A1(n1182), .A2(\completionDataOut[1][15] ), .B1(n1196), 
        .B2(\completionDataOut[3][15] ), .ZN(n1887) );
  AOI22D1 U1749 ( .A1(n1157), .A2(\completionDataOut[0][15] ), .B1(n1170), 
        .B2(\completionDataOut[2][15] ), .ZN(n1886) );
  AOI22D1 U1750 ( .A1(n1179), .A2(\completionDataOut[1][14] ), .B1(n1195), 
        .B2(\completionDataOut[3][14] ), .ZN(n1883) );
  AOI22D1 U1751 ( .A1(n1154), .A2(\completionDataOut[0][14] ), .B1(n1169), 
        .B2(\completionDataOut[2][14] ), .ZN(n1882) );
  AOI22D1 U1752 ( .A1(n1230), .A2(\completionDataOut[5][13] ), .B1(n1245), 
        .B2(\completionDataOut[7][13] ), .ZN(n1881) );
  AOI22D1 U1753 ( .A1(n1205), .A2(\completionDataOut[4][13] ), .B1(n1220), 
        .B2(\completionDataOut[6][13] ), .ZN(n1880) );
  AOI22D1 U1754 ( .A1(n1179), .A2(\completionDataOut[1][13] ), .B1(n1195), 
        .B2(\completionDataOut[3][13] ), .ZN(n1879) );
  AOI22D1 U1755 ( .A1(n1154), .A2(\completionDataOut[0][13] ), .B1(n1169), 
        .B2(\completionDataOut[2][13] ), .ZN(n1878) );
  AOI22D1 U1756 ( .A1(n1230), .A2(\completionDataOut[5][12] ), .B1(n1245), 
        .B2(\completionDataOut[7][12] ), .ZN(n1877) );
  AOI22D1 U1757 ( .A1(n1205), .A2(\completionDataOut[4][12] ), .B1(n1220), 
        .B2(\completionDataOut[6][12] ), .ZN(n1876) );
  AOI22D1 U1758 ( .A1(n1179), .A2(\completionDataOut[1][12] ), .B1(n1195), 
        .B2(\completionDataOut[3][12] ), .ZN(n1875) );
  AOI22D1 U1759 ( .A1(n1154), .A2(\completionDataOut[0][12] ), .B1(n1169), 
        .B2(\completionDataOut[2][12] ), .ZN(n1874) );
  AOI22D1 U1760 ( .A1(n1154), .A2(\completionDataOut[0][11] ), .B1(n1169), 
        .B2(\completionDataOut[2][11] ), .ZN(n1872) );
  AOI22D1 U1761 ( .A1(n1178), .A2(\completionDataOut[1][10] ), .B1(n1190), 
        .B2(\completionDataOut[3][10] ), .ZN(n1869) );
  AOI22D1 U1762 ( .A1(n1153), .A2(\completionDataOut[0][10] ), .B1(n1164), 
        .B2(\completionDataOut[2][10] ), .ZN(n1868) );
  AOI22D1 U1763 ( .A1(n1229), .A2(\completionDataOut[5][9] ), .B1(n1240), .B2(
        \completionDataOut[7][9] ), .ZN(n1867) );
  AOI22D1 U1764 ( .A1(n1204), .A2(\completionDataOut[4][9] ), .B1(n1215), .B2(
        \completionDataOut[6][9] ), .ZN(n1866) );
  AOI22D1 U1765 ( .A1(n1178), .A2(\completionDataOut[1][9] ), .B1(n1190), .B2(
        \completionDataOut[3][9] ), .ZN(n1865) );
  AOI22D1 U1766 ( .A1(n1153), .A2(\completionDataOut[0][9] ), .B1(n1164), .B2(
        \completionDataOut[2][9] ), .ZN(n1864) );
  AOI22D1 U1767 ( .A1(n1153), .A2(\completionDataOut[0][8] ), .B1(n1164), .B2(
        \completionDataOut[2][8] ), .ZN(n1863) );
  AOI22D1 U1768 ( .A1(n1229), .A2(\completionDataOut[5][7] ), .B1(n1240), .B2(
        \completionDataOut[7][7] ), .ZN(n1862) );
  AOI22D1 U1769 ( .A1(n1204), .A2(\completionDataOut[4][7] ), .B1(n1215), .B2(
        \completionDataOut[6][7] ), .ZN(n1861) );
  AOI22D1 U1770 ( .A1(n1178), .A2(\completionDataOut[1][7] ), .B1(n1190), .B2(
        \completionDataOut[3][7] ), .ZN(n1860) );
  AOI22D1 U1771 ( .A1(n1153), .A2(\completionDataOut[0][7] ), .B1(n1164), .B2(
        \completionDataOut[2][7] ), .ZN(n1859) );
  AOI22D1 U1772 ( .A1(n1229), .A2(\completionDataOut[5][6] ), .B1(n1240), .B2(
        \completionDataOut[7][6] ), .ZN(n1858) );
  AOI22D1 U1773 ( .A1(n1178), .A2(\completionDataOut[1][6] ), .B1(n1190), .B2(
        \completionDataOut[3][6] ), .ZN(n1856) );
  AOI22D1 U1774 ( .A1(n1153), .A2(\completionDataOut[0][6] ), .B1(n1164), .B2(
        \completionDataOut[2][6] ), .ZN(n1855) );
  AOI22D1 U1775 ( .A1(n1228), .A2(\completionDataOut[5][5] ), .B1(n1240), .B2(
        \completionDataOut[7][5] ), .ZN(n1854) );
  AOI22D1 U1776 ( .A1(n1203), .A2(\completionDataOut[4][5] ), .B1(n1215), .B2(
        \completionDataOut[6][5] ), .ZN(n1853) );
  AOI22D1 U1777 ( .A1(n1177), .A2(\completionDataOut[1][5] ), .B1(n1190), .B2(
        \completionDataOut[3][5] ), .ZN(n1852) );
  AOI22D1 U1778 ( .A1(n1152), .A2(\completionDataOut[0][5] ), .B1(n1164), .B2(
        \completionDataOut[2][5] ), .ZN(n1851) );
  CKBD1 U1779 ( .I(n1170), .Z(n1164) );
  AOI22D1 U1780 ( .A1(n1228), .A2(\completionDataOut[5][4] ), .B1(n1241), .B2(
        \completionDataOut[7][4] ), .ZN(n1850) );
  AOI22D1 U1781 ( .A1(n1203), .A2(\completionDataOut[4][4] ), .B1(n1216), .B2(
        \completionDataOut[6][4] ), .ZN(n1849) );
  AOI22D1 U1782 ( .A1(n1177), .A2(\completionDataOut[1][4] ), .B1(n1191), .B2(
        \completionDataOut[3][4] ), .ZN(n1848) );
  AOI22D1 U1783 ( .A1(n1152), .A2(\completionDataOut[0][4] ), .B1(n1165), .B2(
        \completionDataOut[2][4] ), .ZN(n1847) );
  AOI22D1 U1784 ( .A1(n1177), .A2(\completionDataOut[1][3] ), .B1(n1191), .B2(
        \completionDataOut[3][3] ), .ZN(n1846) );
  AOI22D1 U1785 ( .A1(n1152), .A2(\completionDataOut[0][3] ), .B1(n1165), .B2(
        \completionDataOut[2][3] ), .ZN(n1845) );
  AOI22D1 U1786 ( .A1(n1152), .A2(\completionDataOut[0][2] ), .B1(n1165), .B2(
        \completionDataOut[2][2] ), .ZN(n1844) );
  AOI22D1 U1787 ( .A1(n1228), .A2(\completionDataOut[5][1] ), .B1(n1241), .B2(
        \completionDataOut[7][1] ), .ZN(n1843) );
  AOI22D1 U1788 ( .A1(n1203), .A2(\completionDataOut[4][1] ), .B1(n1216), .B2(
        \completionDataOut[6][1] ), .ZN(n1842) );
  AOI22D1 U1789 ( .A1(n1177), .A2(\completionDataOut[1][1] ), .B1(n1191), .B2(
        \completionDataOut[3][1] ), .ZN(n1841) );
  AOI22D1 U1790 ( .A1(n1152), .A2(\completionDataOut[0][1] ), .B1(n1165), .B2(
        \completionDataOut[2][1] ), .ZN(n1840) );
  AOI22D1 U1791 ( .A1(n1228), .A2(\completionDataOut[5][0] ), .B1(n1241), .B2(
        \completionDataOut[7][0] ), .ZN(n1839) );
  CKBD1 U1792 ( .I(n1233), .Z(n1229) );
  AOI22D1 U1793 ( .A1(n1203), .A2(\completionDataOut[4][0] ), .B1(n1216), .B2(
        \completionDataOut[6][0] ), .ZN(n1838) );
  CKBD1 U1794 ( .I(n1208), .Z(n1204) );
  AOI22D1 U1795 ( .A1(n1177), .A2(\completionDataOut[1][0] ), .B1(n1191), .B2(
        \completionDataOut[3][0] ), .ZN(n1837) );
  CKBD1 U1796 ( .I(n1182), .Z(n1178) );
  AOI22D1 U1797 ( .A1(n1152), .A2(\completionDataOut[0][0] ), .B1(n1165), .B2(
        \completionDataOut[2][0] ), .ZN(n1836) );
  CKBD1 U1798 ( .I(n1153), .Z(n1152) );
  CKBD1 U1799 ( .I(n1157), .Z(n1153) );
  AOI22D1 U1800 ( .A1(n1026), .A2(\managementDataOut[5][8] ), .B1(n1036), .B2(
        \managementDataOut[7][8] ), .ZN(n1319) );
  AOI22D1 U1801 ( .A1(n994), .A2(\managementDataOut[4][8] ), .B1(n1004), .B2(
        \managementDataOut[6][8] ), .ZN(n1318) );
  AOI22D1 U1802 ( .A1(n964), .A2(\managementDataOut[1][8] ), .B1(n972), .B2(
        \managementDataOut[3][8] ), .ZN(n1317) );
  AOI22D1 U1803 ( .A1(n290), .A2(\managementDataOut[0][8] ), .B1(n954), .B2(
        \managementDataOut[2][8] ), .ZN(n1316) );
  AOI22D1 U1804 ( .A1(n1019), .A2(\managementDataOut[5][7] ), .B1(n1036), .B2(
        \managementDataOut[7][7] ), .ZN(n1323) );
  AOI22D1 U1805 ( .A1(n987), .A2(\managementDataOut[4][7] ), .B1(n1004), .B2(
        \managementDataOut[6][7] ), .ZN(n1322) );
  AOI22D1 U1806 ( .A1(n964), .A2(\managementDataOut[1][7] ), .B1(n972), .B2(
        \managementDataOut[3][7] ), .ZN(n1321) );
  AOI22D1 U1807 ( .A1(n290), .A2(\managementDataOut[0][7] ), .B1(n954), .B2(
        \managementDataOut[2][7] ), .ZN(n1320) );
  AOI22D1 U1808 ( .A1(n1019), .A2(\managementDataOut[5][6] ), .B1(n1036), .B2(
        \managementDataOut[7][6] ), .ZN(n1327) );
  AOI22D1 U1809 ( .A1(n987), .A2(\managementDataOut[4][6] ), .B1(n1004), .B2(
        \managementDataOut[6][6] ), .ZN(n1326) );
  AOI22D1 U1810 ( .A1(n282), .A2(\managementDataOut[1][6] ), .B1(n972), .B2(
        \managementDataOut[3][6] ), .ZN(n1325) );
  AOI22D1 U1811 ( .A1(n286), .A2(\managementDataOut[0][6] ), .B1(n954), .B2(
        \managementDataOut[2][6] ), .ZN(n1324) );
  AOI22D1 U1812 ( .A1(n1019), .A2(\managementDataOut[5][5] ), .B1(n1036), .B2(
        \managementDataOut[7][5] ), .ZN(n1331) );
  AOI22D1 U1813 ( .A1(n987), .A2(\managementDataOut[4][5] ), .B1(n1004), .B2(
        \managementDataOut[6][5] ), .ZN(n1330) );
  AOI22D1 U1814 ( .A1(n274), .A2(\managementDataOut[1][5] ), .B1(n972), .B2(
        \managementDataOut[3][5] ), .ZN(n1329) );
  AOI22D1 U1815 ( .A1(n288), .A2(\managementDataOut[0][5] ), .B1(n954), .B2(
        \managementDataOut[2][5] ), .ZN(n1328) );
  AOI22D1 U1816 ( .A1(n996), .A2(\managementDataOut[4][4] ), .B1(n1004), .B2(
        \managementDataOut[6][4] ), .ZN(n1334) );
  AOI22D1 U1817 ( .A1(n274), .A2(\managementDataOut[1][4] ), .B1(n972), .B2(
        \managementDataOut[3][4] ), .ZN(n1333) );
  AOI22D1 U1818 ( .A1(n294), .A2(\managementDataOut[0][4] ), .B1(n954), .B2(
        \managementDataOut[2][4] ), .ZN(n1332) );
  AOI22D1 U1819 ( .A1(n1019), .A2(\managementDataOut[5][3] ), .B1(n1044), .B2(
        \managementDataOut[7][3] ), .ZN(n1339) );
  AOI22D1 U1820 ( .A1(n987), .A2(\managementDataOut[4][3] ), .B1(n1012), .B2(
        \managementDataOut[6][3] ), .ZN(n1338) );
  AOI22D1 U1821 ( .A1(n278), .A2(\managementDataOut[1][3] ), .B1(n980), .B2(
        \managementDataOut[3][3] ), .ZN(n1337) );
  AOI22D1 U1822 ( .A1(n294), .A2(\managementDataOut[0][3] ), .B1(n962), .B2(
        \managementDataOut[2][3] ), .ZN(n1336) );
  AOI22D1 U1823 ( .A1(n996), .A2(\managementDataOut[4][2] ), .B1(n1008), .B2(
        \managementDataOut[6][2] ), .ZN(n1342) );
  AOI22D1 U1824 ( .A1(n278), .A2(\managementDataOut[1][2] ), .B1(n976), .B2(
        \managementDataOut[3][2] ), .ZN(n1341) );
  AOI22D1 U1825 ( .A1(n1020), .A2(\managementDataOut[5][1] ), .B1(n1043), .B2(
        \managementDataOut[7][1] ), .ZN(n1347) );
  AOI22D1 U1826 ( .A1(n988), .A2(\managementDataOut[4][1] ), .B1(n1011), .B2(
        \managementDataOut[6][1] ), .ZN(n1346) );
  AOI22D1 U1827 ( .A1(n964), .A2(\managementDataOut[1][1] ), .B1(n979), .B2(
        \managementDataOut[3][1] ), .ZN(n1345) );
  AOI22D1 U1828 ( .A1(n290), .A2(\managementDataOut[0][1] ), .B1(n961), .B2(
        \managementDataOut[2][1] ), .ZN(n1344) );
  AOI22D1 U1829 ( .A1(n988), .A2(\managementDataOut[4][0] ), .B1(n1005), .B2(
        \managementDataOut[6][0] ), .ZN(n1350) );
  AOI22D1 U1830 ( .A1(n282), .A2(\managementDataOut[1][0] ), .B1(n973), .B2(
        \managementDataOut[3][0] ), .ZN(n1349) );
  AOI22D1 U1831 ( .A1(n286), .A2(\managementDataOut[0][0] ), .B1(n955), .B2(
        \managementDataOut[2][0] ), .ZN(n1348) );
  AOI22D1 U1832 ( .A1(n988), .A2(\completionDataOut[4][69] ), .B1(n1005), .B2(
        \completionDataOut[6][69] ), .ZN(n1354) );
  AOI22D1 U1833 ( .A1(n276), .A2(\completionDataOut[1][69] ), .B1(n973), .B2(
        \completionDataOut[3][69] ), .ZN(n1353) );
  AOI22D1 U1834 ( .A1(n287), .A2(\completionDataOut[0][69] ), .B1(n955), .B2(
        \completionDataOut[2][69] ), .ZN(n1352) );
  AOI22D1 U1835 ( .A1(n988), .A2(\completionDataOut[4][68] ), .B1(n1005), .B2(
        \completionDataOut[6][68] ), .ZN(n1358) );
  AOI22D1 U1836 ( .A1(n280), .A2(\completionDataOut[1][68] ), .B1(n973), .B2(
        \completionDataOut[3][68] ), .ZN(n1357) );
  AOI22D1 U1837 ( .A1(n297), .A2(\completionDataOut[0][68] ), .B1(n955), .B2(
        \completionDataOut[2][68] ), .ZN(n1356) );
  AOI22D1 U1838 ( .A1(n1020), .A2(\completionDataOut[5][67] ), .B1(n1037), 
        .B2(\completionDataOut[7][67] ), .ZN(n1363) );
  AOI22D1 U1839 ( .A1(n988), .A2(\completionDataOut[4][67] ), .B1(n1005), .B2(
        \completionDataOut[6][67] ), .ZN(n1362) );
  AOI22D1 U1840 ( .A1(n491), .A2(\completionDataOut[1][67] ), .B1(n973), .B2(
        \completionDataOut[3][67] ), .ZN(n1361) );
  AOI22D1 U1841 ( .A1(n293), .A2(\completionDataOut[0][67] ), .B1(n955), .B2(
        \completionDataOut[2][67] ), .ZN(n1360) );
  AOI22D1 U1842 ( .A1(n994), .A2(\completionDataOut[4][66] ), .B1(n1005), .B2(
        \completionDataOut[6][66] ), .ZN(n1366) );
  AOI22D1 U1843 ( .A1(n282), .A2(\completionDataOut[1][66] ), .B1(n973), .B2(
        \completionDataOut[3][66] ), .ZN(n1365) );
  AOI22D1 U1844 ( .A1(n286), .A2(\completionDataOut[0][66] ), .B1(n955), .B2(
        \completionDataOut[2][66] ), .ZN(n1364) );
  AOI22D1 U1845 ( .A1(n986), .A2(\completionDataOut[4][65] ), .B1(n1003), .B2(
        \completionDataOut[6][65] ), .ZN(n1370) );
  AOI22D1 U1846 ( .A1(n283), .A2(\completionDataOut[1][65] ), .B1(n971), .B2(
        \completionDataOut[3][65] ), .ZN(n1369) );
  AOI22D1 U1847 ( .A1(n289), .A2(\completionDataOut[0][65] ), .B1(n953), .B2(
        \completionDataOut[2][65] ), .ZN(n1368) );
  AOI22D1 U1848 ( .A1(n275), .A2(\completionDataOut[1][64] ), .B1(n971), .B2(
        \completionDataOut[3][64] ), .ZN(n1373) );
  AOI22D1 U1849 ( .A1(n286), .A2(\completionDataOut[0][64] ), .B1(n953), .B2(
        \completionDataOut[2][64] ), .ZN(n1372) );
  AOI22D1 U1850 ( .A1(n296), .A2(\completionDataOut[0][63] ), .B1(n953), .B2(
        \completionDataOut[2][63] ), .ZN(n1376) );
  AOI22D1 U1851 ( .A1(n292), .A2(\completionDataOut[0][62] ), .B1(n953), .B2(
        \completionDataOut[2][62] ), .ZN(n1379) );
  AOI22D1 U1852 ( .A1(n279), .A2(\completionDataOut[1][61] ), .B1(n971), .B2(
        \completionDataOut[3][61] ), .ZN(n1383) );
  AOI22D1 U1853 ( .A1(n288), .A2(\completionDataOut[0][61] ), .B1(n953), .B2(
        \completionDataOut[2][61] ), .ZN(n1382) );
  CKBD1 U1854 ( .I(n1043), .Z(n1037) );
  CKBD1 U1855 ( .I(n1011), .Z(n1005) );
  CKBD1 U1856 ( .I(n987), .Z(n988) );
  AOI22D1 U1857 ( .A1(n281), .A2(\completionDataOut[1][60] ), .B1(n971), .B2(
        \completionDataOut[3][60] ), .ZN(n1385) );
  CKBD1 U1858 ( .I(n979), .Z(n973) );
  AOI22D1 U1859 ( .A1(n293), .A2(\completionDataOut[0][60] ), .B1(n953), .B2(
        \completionDataOut[2][60] ), .ZN(n1384) );
  CKBD1 U1860 ( .I(n955), .Z(n953) );
  CKBD1 U1861 ( .I(n961), .Z(n955) );
  AOI22D1 U1862 ( .A1(n1021), .A2(\completionDataOut[5][59] ), .B1(n1038), 
        .B2(\completionDataOut[7][59] ), .ZN(n1389) );
  AOI22D1 U1863 ( .A1(n989), .A2(\completionDataOut[4][59] ), .B1(n1006), .B2(
        \completionDataOut[6][59] ), .ZN(n1388) );
  AOI22D1 U1864 ( .A1(n280), .A2(\completionDataOut[1][59] ), .B1(n974), .B2(
        \completionDataOut[3][59] ), .ZN(n1387) );
  AOI22D1 U1865 ( .A1(n290), .A2(\completionDataOut[0][59] ), .B1(n956), .B2(
        \completionDataOut[2][59] ), .ZN(n1386) );
  AOI22D1 U1866 ( .A1(n285), .A2(\completionDataOut[1][58] ), .B1(n974), .B2(
        \completionDataOut[3][58] ), .ZN(n1391) );
  AOI22D1 U1867 ( .A1(n295), .A2(\completionDataOut[0][58] ), .B1(n956), .B2(
        \completionDataOut[2][58] ), .ZN(n1390) );
  AOI22D1 U1868 ( .A1(n291), .A2(\completionDataOut[0][57] ), .B1(n956), .B2(
        \completionDataOut[2][57] ), .ZN(n1394) );
  AOI22D1 U1869 ( .A1(n287), .A2(\completionDataOut[0][56] ), .B1(n956), .B2(
        \completionDataOut[2][56] ), .ZN(n1396) );
  AOI22D1 U1870 ( .A1(n277), .A2(\completionDataOut[1][55] ), .B1(n976), .B2(
        \completionDataOut[3][55] ), .ZN(n1399) );
  AOI22D1 U1871 ( .A1(n297), .A2(\completionDataOut[0][55] ), .B1(n958), .B2(
        \completionDataOut[2][55] ), .ZN(n1398) );
  AOI22D1 U1872 ( .A1(n994), .A2(\completionDataOut[4][54] ), .B1(n1008), .B2(
        \completionDataOut[6][54] ), .ZN(n1402) );
  AOI22D1 U1873 ( .A1(n274), .A2(\completionDataOut[1][54] ), .B1(n976), .B2(
        \completionDataOut[3][54] ), .ZN(n1401) );
  AOI22D1 U1874 ( .A1(n289), .A2(\completionDataOut[0][54] ), .B1(n958), .B2(
        \completionDataOut[2][54] ), .ZN(n1400) );
  AOI22D1 U1875 ( .A1(n1227), .A2(\completionDataOut[5][19] ), .B1(n1239), 
        .B2(\completionDataOut[7][19] ), .ZN(n1901) );
  AOI22D1 U1876 ( .A1(n1202), .A2(\completionDataOut[4][19] ), .B1(n1214), 
        .B2(\completionDataOut[6][19] ), .ZN(n1900) );
  AOI22D1 U1877 ( .A1(n1176), .A2(\completionDataOut[1][19] ), .B1(n1189), 
        .B2(\completionDataOut[3][19] ), .ZN(n1899) );
  AOI22D1 U1878 ( .A1(n1151), .A2(\completionDataOut[0][19] ), .B1(n1163), 
        .B2(\completionDataOut[2][19] ), .ZN(n1898) );
  AOI22D1 U1879 ( .A1(n1017), .A2(\completionDataOut[5][53] ), .B1(n1034), 
        .B2(\completionDataOut[7][53] ), .ZN(n1407) );
  AOI22D1 U1880 ( .A1(n985), .A2(\completionDataOut[4][53] ), .B1(n1002), .B2(
        \completionDataOut[6][53] ), .ZN(n1406) );
  AOI22D1 U1881 ( .A1(n278), .A2(\completionDataOut[1][53] ), .B1(n970), .B2(
        \completionDataOut[3][53] ), .ZN(n1405) );
  AOI22D1 U1882 ( .A1(n297), .A2(\completionDataOut[0][53] ), .B1(n952), .B2(
        \completionDataOut[2][53] ), .ZN(n1404) );
  AOI22D1 U1883 ( .A1(n1017), .A2(\completionDataOut[5][52] ), .B1(n1034), 
        .B2(\completionDataOut[7][52] ), .ZN(n1411) );
  AOI22D1 U1884 ( .A1(n985), .A2(\completionDataOut[4][52] ), .B1(n1002), .B2(
        \completionDataOut[6][52] ), .ZN(n1410) );
  AOI22D1 U1885 ( .A1(n280), .A2(\completionDataOut[1][52] ), .B1(n970), .B2(
        \completionDataOut[3][52] ), .ZN(n1409) );
  AOI22D1 U1886 ( .A1(n293), .A2(\completionDataOut[0][52] ), .B1(n952), .B2(
        \completionDataOut[2][52] ), .ZN(n1408) );
  AOI22D1 U1887 ( .A1(n1017), .A2(\completionDataOut[5][51] ), .B1(n1034), 
        .B2(\completionDataOut[7][51] ), .ZN(n1415) );
  AOI22D1 U1888 ( .A1(n985), .A2(\completionDataOut[4][51] ), .B1(n1002), .B2(
        \completionDataOut[6][51] ), .ZN(n1414) );
  AOI22D1 U1889 ( .A1(n276), .A2(\completionDataOut[1][51] ), .B1(n970), .B2(
        \completionDataOut[3][51] ), .ZN(n1413) );
  AOI22D1 U1890 ( .A1(n289), .A2(\completionDataOut[0][51] ), .B1(n952), .B2(
        \completionDataOut[2][51] ), .ZN(n1412) );
  AOI22D1 U1891 ( .A1(n1017), .A2(\completionDataOut[5][50] ), .B1(n1034), 
        .B2(\completionDataOut[7][50] ), .ZN(n1419) );
  AOI22D1 U1892 ( .A1(n985), .A2(\completionDataOut[4][50] ), .B1(n1002), .B2(
        \completionDataOut[6][50] ), .ZN(n1418) );
  AOI22D1 U1893 ( .A1(n281), .A2(\completionDataOut[1][50] ), .B1(n970), .B2(
        \completionDataOut[3][50] ), .ZN(n1417) );
  AOI22D1 U1894 ( .A1(n296), .A2(\completionDataOut[0][50] ), .B1(n952), .B2(
        \completionDataOut[2][50] ), .ZN(n1416) );
  AOI22D1 U1895 ( .A1(n296), .A2(\completionDataOut[0][49] ), .B1(n952), .B2(
        \completionDataOut[2][49] ), .ZN(n1420) );
  CKBD1 U1896 ( .I(n1026), .Z(n1021) );
  AOI22D1 U1897 ( .A1(n284), .A2(\completionDataOut[1][48] ), .B1(n970), .B2(
        \completionDataOut[3][48] ), .ZN(n1423) );
  CKBD1 U1898 ( .I(n974), .Z(n970) );
  AOI22D1 U1899 ( .A1(n292), .A2(\completionDataOut[0][48] ), .B1(n952), .B2(
        \completionDataOut[2][48] ), .ZN(n1422) );
  CKBD1 U1900 ( .I(n956), .Z(n952) );
  AOI22D1 U1901 ( .A1(n990), .A2(\completionDataOut[4][47] ), .B1(n1007), .B2(
        \completionDataOut[6][47] ), .ZN(n1426) );
  AOI22D1 U1902 ( .A1(n285), .A2(\completionDataOut[1][47] ), .B1(n975), .B2(
        \completionDataOut[3][47] ), .ZN(n1425) );
  AOI22D1 U1903 ( .A1(n295), .A2(\completionDataOut[0][47] ), .B1(n957), .B2(
        \completionDataOut[2][47] ), .ZN(n1424) );
  AOI22D1 U1904 ( .A1(n277), .A2(\completionDataOut[1][46] ), .B1(n975), .B2(
        \completionDataOut[3][46] ), .ZN(n1428) );
  AOI22D1 U1905 ( .A1(n291), .A2(\completionDataOut[0][46] ), .B1(n957), .B2(
        \completionDataOut[2][46] ), .ZN(n1427) );
  AOI22D1 U1906 ( .A1(n990), .A2(\completionDataOut[4][45] ), .B1(n1007), .B2(
        \completionDataOut[6][45] ), .ZN(n1433) );
  AOI22D1 U1907 ( .A1(n281), .A2(\completionDataOut[1][45] ), .B1(n975), .B2(
        \completionDataOut[3][45] ), .ZN(n1432) );
  AOI22D1 U1908 ( .A1(n287), .A2(\completionDataOut[0][45] ), .B1(n957), .B2(
        \completionDataOut[2][45] ), .ZN(n1431) );
  AOI22D1 U1909 ( .A1(n285), .A2(\completionDataOut[1][44] ), .B1(n979), .B2(
        \completionDataOut[3][44] ), .ZN(n1436) );
  AOI22D1 U1910 ( .A1(n292), .A2(\completionDataOut[0][44] ), .B1(n961), .B2(
        \completionDataOut[2][44] ), .ZN(n1435) );
  AOI22D1 U1911 ( .A1(n297), .A2(\completionDataOut[0][43] ), .B1(n957), .B2(
        \completionDataOut[2][43] ), .ZN(n1438) );
  AOI22D1 U1912 ( .A1(n278), .A2(\completionDataOut[1][42] ), .B1(n979), .B2(
        \completionDataOut[3][42] ), .ZN(n1440) );
  AOI22D1 U1913 ( .A1(n294), .A2(\completionDataOut[0][42] ), .B1(n961), .B2(
        \completionDataOut[2][42] ), .ZN(n1439) );
  AOI22D1 U1914 ( .A1(n1016), .A2(\completionDataOut[5][41] ), .B1(n1033), 
        .B2(\completionDataOut[7][41] ), .ZN(n1445) );
  AOI22D1 U1915 ( .A1(n984), .A2(\completionDataOut[4][41] ), .B1(n1001), .B2(
        \completionDataOut[6][41] ), .ZN(n1444) );
  AOI22D1 U1916 ( .A1(n276), .A2(\completionDataOut[1][41] ), .B1(n969), .B2(
        \completionDataOut[3][41] ), .ZN(n1443) );
  AOI22D1 U1917 ( .A1(n293), .A2(\completionDataOut[0][41] ), .B1(n951), .B2(
        \completionDataOut[2][41] ), .ZN(n1442) );
  AOI22D1 U1918 ( .A1(n280), .A2(\completionDataOut[1][40] ), .B1(n969), .B2(
        \completionDataOut[3][40] ), .ZN(n1447) );
  AOI22D1 U1919 ( .A1(n289), .A2(\completionDataOut[0][40] ), .B1(n951), .B2(
        \completionDataOut[2][40] ), .ZN(n1446) );
  AOI22D1 U1920 ( .A1(n1016), .A2(\completionDataOut[5][39] ), .B1(n1033), 
        .B2(\completionDataOut[7][39] ), .ZN(n1453) );
  AOI22D1 U1921 ( .A1(n984), .A2(\completionDataOut[4][39] ), .B1(n1001), .B2(
        \completionDataOut[6][39] ), .ZN(n1452) );
  AOI22D1 U1922 ( .A1(n284), .A2(\completionDataOut[1][39] ), .B1(n969), .B2(
        \completionDataOut[3][39] ), .ZN(n1451) );
  AOI22D1 U1923 ( .A1(n291), .A2(\completionDataOut[0][39] ), .B1(n951), .B2(
        \completionDataOut[2][39] ), .ZN(n1450) );
  AOI22D1 U1924 ( .A1(n1016), .A2(\completionDataOut[5][38] ), .B1(n1033), 
        .B2(\completionDataOut[7][38] ), .ZN(n1457) );
  AOI22D1 U1925 ( .A1(n984), .A2(\completionDataOut[4][38] ), .B1(n1001), .B2(
        \completionDataOut[6][38] ), .ZN(n1456) );
  AOI22D1 U1926 ( .A1(n283), .A2(\completionDataOut[1][38] ), .B1(n969), .B2(
        \completionDataOut[3][38] ), .ZN(n1455) );
  AOI22D1 U1927 ( .A1(n296), .A2(\completionDataOut[0][38] ), .B1(n951), .B2(
        \completionDataOut[2][38] ), .ZN(n1454) );
  AOI22D1 U1928 ( .A1(n275), .A2(\completionDataOut[1][36] ), .B1(n969), .B2(
        \completionDataOut[3][36] ), .ZN(n1463) );
  AOI22D1 U1929 ( .A1(n292), .A2(\completionDataOut[0][36] ), .B1(n951), .B2(
        \completionDataOut[2][36] ), .ZN(n1462) );
  AOI22D1 U1930 ( .A1(n1023), .A2(\completionDataOut[5][35] ), .B1(n1032), 
        .B2(\completionDataOut[7][35] ), .ZN(n1467) );
  AOI22D1 U1931 ( .A1(n991), .A2(\completionDataOut[4][35] ), .B1(n1000), .B2(
        \completionDataOut[6][35] ), .ZN(n1466) );
  AOI22D1 U1932 ( .A1(n964), .A2(\completionDataOut[1][35] ), .B1(n968), .B2(
        \completionDataOut[3][35] ), .ZN(n1465) );
  AOI22D1 U1933 ( .A1(n292), .A2(\completionDataOut[0][35] ), .B1(n950), .B2(
        \completionDataOut[2][35] ), .ZN(n1464) );
  AOI22D1 U1934 ( .A1(n283), .A2(\completionDataOut[1][34] ), .B1(n968), .B2(
        \completionDataOut[3][34] ), .ZN(n1469) );
  AOI22D1 U1935 ( .A1(n288), .A2(\completionDataOut[0][34] ), .B1(n950), .B2(
        \completionDataOut[2][34] ), .ZN(n1468) );
  AOI22D1 U1936 ( .A1(n275), .A2(\completionDataOut[1][33] ), .B1(n968), .B2(
        \completionDataOut[3][33] ), .ZN(n1473) );
  AOI22D1 U1937 ( .A1(n945), .A2(\completionDataOut[0][33] ), .B1(n950), .B2(
        \completionDataOut[2][33] ), .ZN(n1472) );
  AOI22D1 U1938 ( .A1(n279), .A2(\completionDataOut[1][32] ), .B1(n968), .B2(
        \completionDataOut[3][32] ), .ZN(n1477) );
  AOI22D1 U1939 ( .A1(n295), .A2(\completionDataOut[0][32] ), .B1(n950), .B2(
        \completionDataOut[2][32] ), .ZN(n1476) );
  AOI22D1 U1940 ( .A1(n291), .A2(\completionDataOut[0][31] ), .B1(n950), .B2(
        \completionDataOut[2][31] ), .ZN(n1480) );
  AOI22D1 U1941 ( .A1(n1025), .A2(\completionDataOut[5][30] ), .B1(n1032), 
        .B2(\completionDataOut[7][30] ), .ZN(n1485) );
  CKBD1 U1942 ( .I(n1040), .Z(n1032) );
  AOI22D1 U1943 ( .A1(n993), .A2(\completionDataOut[4][30] ), .B1(n1000), .B2(
        \completionDataOut[6][30] ), .ZN(n1484) );
  CKBD1 U1944 ( .I(n1008), .Z(n1000) );
  AOI22D1 U1945 ( .A1(n491), .A2(\completionDataOut[1][30] ), .B1(n968), .B2(
        \completionDataOut[3][30] ), .ZN(n1483) );
  CKBD1 U1946 ( .I(n976), .Z(n968) );
  AOI22D1 U1947 ( .A1(n286), .A2(\completionDataOut[0][30] ), .B1(n950), .B2(
        \completionDataOut[2][30] ), .ZN(n1482) );
  CKBD1 U1948 ( .I(n958), .Z(n950) );
  AOI22D1 U1949 ( .A1(n1015), .A2(\completionDataOut[5][29] ), .B1(n1031), 
        .B2(\completionDataOut[7][29] ), .ZN(n1489) );
  AOI22D1 U1950 ( .A1(n983), .A2(\completionDataOut[4][29] ), .B1(n999), .B2(
        \completionDataOut[6][29] ), .ZN(n1488) );
  AOI22D1 U1951 ( .A1(n285), .A2(\completionDataOut[1][29] ), .B1(n967), .B2(
        \completionDataOut[3][29] ), .ZN(n1487) );
  AOI22D1 U1952 ( .A1(n287), .A2(\completionDataOut[0][29] ), .B1(n949), .B2(
        \completionDataOut[2][29] ), .ZN(n1486) );
  AOI22D1 U1953 ( .A1(n1015), .A2(\completionDataOut[5][28] ), .B1(n1031), 
        .B2(\completionDataOut[7][28] ), .ZN(n1493) );
  AOI22D1 U1954 ( .A1(n983), .A2(\completionDataOut[4][28] ), .B1(n999), .B2(
        \completionDataOut[6][28] ), .ZN(n1492) );
  AOI22D1 U1955 ( .A1(n277), .A2(\completionDataOut[1][28] ), .B1(n967), .B2(
        \completionDataOut[3][28] ), .ZN(n1491) );
  AOI22D1 U1956 ( .A1(n945), .A2(\completionDataOut[0][28] ), .B1(n949), .B2(
        \completionDataOut[2][28] ), .ZN(n1490) );
  AOI22D1 U1957 ( .A1(n281), .A2(\completionDataOut[1][27] ), .B1(n967), .B2(
        \completionDataOut[3][27] ), .ZN(n1495) );
  AOI22D1 U1958 ( .A1(n297), .A2(\completionDataOut[0][27] ), .B1(n949), .B2(
        \completionDataOut[2][27] ), .ZN(n1494) );
  AOI22D1 U1959 ( .A1(n963), .A2(\completionDataOut[1][26] ), .B1(n967), .B2(
        \completionDataOut[3][26] ), .ZN(n1499) );
  AOI22D1 U1960 ( .A1(n293), .A2(\completionDataOut[0][26] ), .B1(n949), .B2(
        \completionDataOut[2][26] ), .ZN(n1498) );
  AOI22D1 U1961 ( .A1(n1015), .A2(\completionDataOut[5][25] ), .B1(n1031), 
        .B2(\completionDataOut[7][25] ), .ZN(n1505) );
  AOI22D1 U1962 ( .A1(n983), .A2(\completionDataOut[4][25] ), .B1(n999), .B2(
        \completionDataOut[6][25] ), .ZN(n1504) );
  AOI22D1 U1963 ( .A1(n284), .A2(\completionDataOut[1][25] ), .B1(n967), .B2(
        \completionDataOut[3][25] ), .ZN(n1503) );
  AOI22D1 U1964 ( .A1(n289), .A2(\completionDataOut[0][25] ), .B1(n949), .B2(
        \completionDataOut[2][25] ), .ZN(n1502) );
  CKBD1 U1965 ( .I(n1040), .Z(n1031) );
  CKBD1 U1966 ( .I(n1044), .Z(n1036) );
  CKBD1 U1967 ( .I(n1025), .Z(n1023) );
  CKBD1 U1968 ( .I(n1008), .Z(n999) );
  CKBD1 U1969 ( .I(n1012), .Z(n1004) );
  CKBD1 U1970 ( .I(n993), .Z(n991) );
  AOI22D1 U1971 ( .A1(n276), .A2(\completionDataOut[1][24] ), .B1(n967), .B2(
        \completionDataOut[3][24] ), .ZN(n1507) );
  CKBD1 U1972 ( .I(n976), .Z(n967) );
  CKBD1 U1973 ( .I(n972), .Z(n976) );
  CKBD1 U1974 ( .I(n980), .Z(n972) );
  AOI22D1 U1975 ( .A1(n945), .A2(\completionDataOut[0][24] ), .B1(n949), .B2(
        \completionDataOut[2][24] ), .ZN(n1506) );
  CKBD1 U1976 ( .I(n958), .Z(n949) );
  CKBD1 U1977 ( .I(n954), .Z(n958) );
  CKBD1 U1978 ( .I(n962), .Z(n954) );
  AOI22D1 U1979 ( .A1(n1027), .A2(\completionDataOut[5][23] ), .B1(n1041), 
        .B2(\completionDataOut[7][23] ), .ZN(n1511) );
  AOI22D1 U1980 ( .A1(n995), .A2(\completionDataOut[4][23] ), .B1(n1009), .B2(
        \completionDataOut[6][23] ), .ZN(n1510) );
  AOI22D1 U1981 ( .A1(n282), .A2(\completionDataOut[1][23] ), .B1(n977), .B2(
        \completionDataOut[3][23] ), .ZN(n1509) );
  AOI22D1 U1982 ( .A1(n945), .A2(\completionDataOut[0][23] ), .B1(n959), .B2(
        \completionDataOut[2][23] ), .ZN(n1508) );
  AOI22D1 U1983 ( .A1(n964), .A2(\completionDataOut[1][22] ), .B1(n977), .B2(
        \completionDataOut[3][22] ), .ZN(n1513) );
  AOI22D1 U1984 ( .A1(n286), .A2(\completionDataOut[0][22] ), .B1(n959), .B2(
        \completionDataOut[2][22] ), .ZN(n1512) );
  AOI22D1 U1985 ( .A1(n278), .A2(\completionDataOut[1][21] ), .B1(n977), .B2(
        \completionDataOut[3][21] ), .ZN(n1517) );
  AOI22D1 U1986 ( .A1(n290), .A2(\completionDataOut[0][21] ), .B1(n959), .B2(
        \completionDataOut[2][21] ), .ZN(n1516) );
  AOI22D1 U1987 ( .A1(n274), .A2(\completionDataOut[1][20] ), .B1(n977), .B2(
        \completionDataOut[3][20] ), .ZN(n1521) );
  AOI22D1 U1988 ( .A1(n294), .A2(\completionDataOut[0][20] ), .B1(n959), .B2(
        \completionDataOut[2][20] ), .ZN(n1520) );
  AOI22D1 U1989 ( .A1(n946), .A2(\completionDataOut[0][19] ), .B1(n959), .B2(
        \completionDataOut[2][19] ), .ZN(n1524) );
  AOI22D1 U1990 ( .A1(n1025), .A2(\completionDataOut[5][18] ), .B1(n1044), 
        .B2(\completionDataOut[7][18] ), .ZN(n1527) );
  AOI22D1 U1991 ( .A1(n278), .A2(\completionDataOut[1][18] ), .B1(n980), .B2(
        \completionDataOut[3][18] ), .ZN(n1526) );
  AOI22D1 U1992 ( .A1(n290), .A2(\completionDataOut[0][18] ), .B1(n962), .B2(
        \completionDataOut[2][18] ), .ZN(n1525) );
  AOI22D1 U1993 ( .A1(n1014), .A2(\completionDataOut[5][17] ), .B1(n1030), 
        .B2(\completionDataOut[7][17] ), .ZN(n1531) );
  AOI22D1 U1994 ( .A1(n982), .A2(\completionDataOut[4][17] ), .B1(n998), .B2(
        \completionDataOut[6][17] ), .ZN(n1530) );
  AOI22D1 U1995 ( .A1(n280), .A2(\completionDataOut[1][17] ), .B1(n966), .B2(
        \completionDataOut[3][17] ), .ZN(n1529) );
  AOI22D1 U1996 ( .A1(n296), .A2(\completionDataOut[0][17] ), .B1(n948), .B2(
        \completionDataOut[2][17] ), .ZN(n1528) );
  AOI22D1 U1997 ( .A1(n963), .A2(\completionDataOut[1][16] ), .B1(n966), .B2(
        \completionDataOut[3][16] ), .ZN(n1533) );
  AOI22D1 U1998 ( .A1(n292), .A2(\completionDataOut[0][16] ), .B1(n948), .B2(
        \completionDataOut[2][16] ), .ZN(n1532) );
  AOI22D1 U1999 ( .A1(n1014), .A2(\completionDataOut[5][15] ), .B1(n1030), 
        .B2(\completionDataOut[7][15] ), .ZN(n1539) );
  AOI22D1 U2000 ( .A1(n982), .A2(\completionDataOut[4][15] ), .B1(n998), .B2(
        \completionDataOut[6][15] ), .ZN(n1538) );
  AOI22D1 U2001 ( .A1(n283), .A2(\completionDataOut[1][15] ), .B1(n966), .B2(
        \completionDataOut[3][15] ), .ZN(n1537) );
  AOI22D1 U2002 ( .A1(n288), .A2(\completionDataOut[0][15] ), .B1(n948), .B2(
        \completionDataOut[2][15] ), .ZN(n1536) );
  AOI22D1 U2003 ( .A1(n275), .A2(\completionDataOut[1][14] ), .B1(n966), .B2(
        \completionDataOut[3][14] ), .ZN(n1541) );
  AOI22D1 U2004 ( .A1(n295), .A2(\completionDataOut[0][14] ), .B1(n948), .B2(
        \completionDataOut[2][14] ), .ZN(n1540) );
  AOI22D1 U2005 ( .A1(n1014), .A2(\completionDataOut[5][13] ), .B1(n1030), 
        .B2(\completionDataOut[7][13] ), .ZN(n1547) );
  AOI22D1 U2006 ( .A1(n982), .A2(\completionDataOut[4][13] ), .B1(n998), .B2(
        \completionDataOut[6][13] ), .ZN(n1546) );
  AOI22D1 U2007 ( .A1(n279), .A2(\completionDataOut[1][13] ), .B1(n966), .B2(
        \completionDataOut[3][13] ), .ZN(n1545) );
  AOI22D1 U2008 ( .A1(n291), .A2(\completionDataOut[0][13] ), .B1(n948), .B2(
        \completionDataOut[2][13] ), .ZN(n1544) );
  CKBD1 U2009 ( .I(n1044), .Z(n1041) );
  CKBD1 U2010 ( .I(n1025), .Z(n1014) );
  CKBD1 U2011 ( .I(n1012), .Z(n1009) );
  AOI22D1 U2012 ( .A1(n287), .A2(\completionDataOut[0][12] ), .B1(n948), .B2(
        \completionDataOut[2][12] ), .ZN(n1548) );
  CKBD1 U2013 ( .I(n959), .Z(n948) );
  CKBD1 U2014 ( .I(n962), .Z(n959) );
  AOI22D1 U2015 ( .A1(n1024), .A2(\completionDataOut[5][11] ), .B1(n1042), 
        .B2(\completionDataOut[7][11] ), .ZN(n1553) );
  AOI22D1 U2016 ( .A1(n992), .A2(\completionDataOut[4][11] ), .B1(n1010), .B2(
        \completionDataOut[6][11] ), .ZN(n1552) );
  AOI22D1 U2017 ( .A1(n283), .A2(\completionDataOut[1][11] ), .B1(n978), .B2(
        \completionDataOut[3][11] ), .ZN(n1551) );
  AOI22D1 U2018 ( .A1(n288), .A2(\completionDataOut[0][11] ), .B1(n960), .B2(
        \completionDataOut[2][11] ), .ZN(n1550) );
  AOI22D1 U2019 ( .A1(n275), .A2(\completionDataOut[1][10] ), .B1(n978), .B2(
        \completionDataOut[3][10] ), .ZN(n1555) );
  AOI22D1 U2020 ( .A1(n295), .A2(\completionDataOut[0][10] ), .B1(n960), .B2(
        \completionDataOut[2][10] ), .ZN(n1554) );
  AOI22D1 U2021 ( .A1(n1024), .A2(\completionDataOut[5][9] ), .B1(n1042), .B2(
        \completionDataOut[7][9] ), .ZN(n1561) );
  AOI22D1 U2022 ( .A1(n992), .A2(\completionDataOut[4][9] ), .B1(n1010), .B2(
        \completionDataOut[6][9] ), .ZN(n1560) );
  AOI22D1 U2023 ( .A1(n279), .A2(\completionDataOut[1][9] ), .B1(n978), .B2(
        \completionDataOut[3][9] ), .ZN(n1559) );
  AOI22D1 U2024 ( .A1(n295), .A2(\completionDataOut[0][9] ), .B1(n960), .B2(
        \completionDataOut[2][9] ), .ZN(n1558) );
  AOI22D1 U2025 ( .A1(n1024), .A2(\completionDataOut[5][8] ), .B1(n1042), .B2(
        \completionDataOut[7][8] ), .ZN(n1565) );
  AOI22D1 U2026 ( .A1(n992), .A2(\completionDataOut[4][8] ), .B1(n1010), .B2(
        \completionDataOut[6][8] ), .ZN(n1564) );
  AOI22D1 U2027 ( .A1(n283), .A2(\completionDataOut[1][8] ), .B1(n978), .B2(
        \completionDataOut[3][8] ), .ZN(n1563) );
  AOI22D1 U2028 ( .A1(n291), .A2(\completionDataOut[0][8] ), .B1(n960), .B2(
        \completionDataOut[2][8] ), .ZN(n1562) );
  AOI22D1 U2029 ( .A1(n287), .A2(\completionDataOut[0][7] ), .B1(n960), .B2(
        \completionDataOut[2][7] ), .ZN(n1566) );
  AOI22D1 U2030 ( .A1(n274), .A2(\completionDataOut[1][6] ), .B1(n980), .B2(
        \completionDataOut[3][6] ), .ZN(n1568) );
  AOI22D1 U2031 ( .A1(n294), .A2(\completionDataOut[0][6] ), .B1(n962), .B2(
        \completionDataOut[2][6] ), .ZN(n1567) );
  AOI22D1 U2032 ( .A1(n1013), .A2(\completionDataOut[5][5] ), .B1(n1029), .B2(
        \completionDataOut[7][5] ), .ZN(n1573) );
  AOI22D1 U2033 ( .A1(n981), .A2(\completionDataOut[4][5] ), .B1(n997), .B2(
        \completionDataOut[6][5] ), .ZN(n1572) );
  AOI22D1 U2034 ( .A1(n277), .A2(\completionDataOut[1][5] ), .B1(n965), .B2(
        \completionDataOut[3][5] ), .ZN(n1571) );
  AOI22D1 U2035 ( .A1(n294), .A2(\completionDataOut[0][5] ), .B1(n947), .B2(
        \completionDataOut[2][5] ), .ZN(n1570) );
  AOI22D1 U2036 ( .A1(n1013), .A2(\completionDataOut[5][4] ), .B1(n1029), .B2(
        \completionDataOut[7][4] ), .ZN(n1577) );
  AOI22D1 U2037 ( .A1(n981), .A2(\completionDataOut[4][4] ), .B1(n997), .B2(
        \completionDataOut[6][4] ), .ZN(n1576) );
  AOI22D1 U2038 ( .A1(n281), .A2(\completionDataOut[1][4] ), .B1(n965), .B2(
        \completionDataOut[3][4] ), .ZN(n1575) );
  AOI22D1 U2039 ( .A1(n297), .A2(\completionDataOut[0][4] ), .B1(n947), .B2(
        \completionDataOut[2][4] ), .ZN(n1574) );
  AOI22D1 U2040 ( .A1(n1013), .A2(\completionDataOut[5][3] ), .B1(n1029), .B2(
        \completionDataOut[7][3] ), .ZN(n1581) );
  AOI22D1 U2041 ( .A1(n981), .A2(\completionDataOut[4][3] ), .B1(n997), .B2(
        \completionDataOut[6][3] ), .ZN(n1580) );
  AOI22D1 U2042 ( .A1(n282), .A2(\completionDataOut[1][3] ), .B1(n965), .B2(
        \completionDataOut[3][3] ), .ZN(n1579) );
  AOI22D1 U2043 ( .A1(n293), .A2(\completionDataOut[0][3] ), .B1(n947), .B2(
        \completionDataOut[2][3] ), .ZN(n1578) );
  AOI22D1 U2044 ( .A1(n1013), .A2(\completionDataOut[5][2] ), .B1(n1029), .B2(
        \completionDataOut[7][2] ), .ZN(n1585) );
  AOI22D1 U2045 ( .A1(n981), .A2(\completionDataOut[4][2] ), .B1(n997), .B2(
        \completionDataOut[6][2] ), .ZN(n1584) );
  AOI22D1 U2046 ( .A1(n284), .A2(\completionDataOut[1][2] ), .B1(n965), .B2(
        \completionDataOut[3][2] ), .ZN(n1583) );
  AOI22D1 U2047 ( .A1(n289), .A2(\completionDataOut[0][2] ), .B1(n947), .B2(
        \completionDataOut[2][2] ), .ZN(n1582) );
  AOI22D1 U2048 ( .A1(n276), .A2(\completionDataOut[1][1] ), .B1(n965), .B2(
        \completionDataOut[3][1] ), .ZN(n1587) );
  AOI22D1 U2049 ( .A1(n946), .A2(\completionDataOut[0][1] ), .B1(n947), .B2(
        \completionDataOut[2][1] ), .ZN(n1586) );
  CKBD1 U2050 ( .I(n1044), .Z(n1042) );
  CKBD1 U2051 ( .I(n1043), .Z(n1038) );
  CKBD1 U2052 ( .I(n1025), .Z(n1024) );
  CKBD1 U2053 ( .I(n1028), .Z(n1027) );
  CKBD1 U2054 ( .I(n1011), .Z(n1006) );
  CKBD1 U2055 ( .I(n996), .Z(n995) );
  CKBD1 U2056 ( .I(n978), .Z(n965) );
  AOI22D1 U2057 ( .A1(n296), .A2(\completionDataOut[0][0] ), .B1(n947), .B2(
        \completionDataOut[2][0] ), .ZN(n1588) );
  CKBD1 U2058 ( .I(n960), .Z(n947) );
  CKBD1 U2059 ( .I(n962), .Z(n960) );
  CKBD1 U2060 ( .I(n961), .Z(n956) );
  AOI22D1 U2061 ( .A1(n1176), .A2(\completionDataOut[1][20] ), .B1(n1189), 
        .B2(\completionDataOut[3][20] ), .ZN(n1903) );
  AOI22D1 U2062 ( .A1(n1151), .A2(\completionDataOut[0][20] ), .B1(n1163), 
        .B2(\completionDataOut[2][20] ), .ZN(n1902) );
  AOI22D1 U2063 ( .A1(n1106), .A2(\completionDataOut[4][61] ), .B1(n1108), 
        .B2(\completionDataOut[6][61] ), .ZN(n1812) );
  AOI22D1 U2064 ( .A1(n1130), .A2(\completionDataOut[5][60] ), .B1(n1133), 
        .B2(\completionDataOut[7][60] ), .ZN(n1811) );
  AOI22D1 U2065 ( .A1(n1106), .A2(\completionDataOut[4][60] ), .B1(n1108), 
        .B2(\completionDataOut[6][60] ), .ZN(n1810) );
  AOI22D1 U2066 ( .A1(n1080), .A2(\completionDataOut[1][60] ), .B1(n1083), 
        .B2(\completionDataOut[3][60] ), .ZN(n1809) );
  AOI22D1 U2067 ( .A1(n1055), .A2(\completionDataOut[0][60] ), .B1(n1057), 
        .B2(\completionDataOut[2][60] ), .ZN(n1808) );
  AOI22D1 U2068 ( .A1(n1130), .A2(\completionDataOut[5][59] ), .B1(n1133), 
        .B2(\completionDataOut[7][59] ), .ZN(n1807) );
  AOI22D1 U2069 ( .A1(n1106), .A2(\completionDataOut[4][59] ), .B1(n1108), 
        .B2(\completionDataOut[6][59] ), .ZN(n1806) );
  AOI22D1 U2070 ( .A1(n1080), .A2(\completionDataOut[1][59] ), .B1(n1083), 
        .B2(\completionDataOut[3][59] ), .ZN(n1805) );
  AOI22D1 U2071 ( .A1(n1055), .A2(\completionDataOut[0][59] ), .B1(n1057), 
        .B2(\completionDataOut[2][59] ), .ZN(n1804) );
  AOI22D1 U2072 ( .A1(n1070), .A2(\completionDataOut[1][58] ), .B1(n1084), 
        .B2(\completionDataOut[3][58] ), .ZN(n1801) );
  AOI22D1 U2073 ( .A1(n1045), .A2(\completionDataOut[0][58] ), .B1(n1058), 
        .B2(\completionDataOut[2][58] ), .ZN(n1800) );
  AOI22D1 U2074 ( .A1(n1096), .A2(\completionDataOut[4][57] ), .B1(n1109), 
        .B2(\completionDataOut[6][57] ), .ZN(n1798) );
  AOI22D1 U2075 ( .A1(n1070), .A2(\completionDataOut[1][57] ), .B1(n1084), 
        .B2(\completionDataOut[3][57] ), .ZN(n1797) );
  AOI22D1 U2076 ( .A1(n1045), .A2(\completionDataOut[0][57] ), .B1(n1058), 
        .B2(\completionDataOut[2][57] ), .ZN(n1796) );
  AOI22D1 U2077 ( .A1(n1096), .A2(\completionDataOut[4][56] ), .B1(n1109), 
        .B2(\completionDataOut[6][56] ), .ZN(n1794) );
  AOI22D1 U2078 ( .A1(n1070), .A2(\completionDataOut[1][56] ), .B1(n1084), 
        .B2(\completionDataOut[3][56] ), .ZN(n1793) );
  AOI22D1 U2079 ( .A1(n1045), .A2(\completionDataOut[0][56] ), .B1(n1058), 
        .B2(\completionDataOut[2][56] ), .ZN(n1792) );
  AOI22D1 U2080 ( .A1(n1120), .A2(\completionDataOut[5][55] ), .B1(n1134), 
        .B2(\completionDataOut[7][55] ), .ZN(n1791) );
  AOI22D1 U2081 ( .A1(n1096), .A2(\completionDataOut[4][55] ), .B1(n1109), 
        .B2(\completionDataOut[6][55] ), .ZN(n1790) );
  AOI22D1 U2082 ( .A1(n1070), .A2(\completionDataOut[1][55] ), .B1(n1084), 
        .B2(\completionDataOut[3][55] ), .ZN(n1789) );
  AOI22D1 U2083 ( .A1(n1045), .A2(\completionDataOut[0][55] ), .B1(n1058), 
        .B2(\completionDataOut[2][55] ), .ZN(n1788) );
  AOI22D1 U2084 ( .A1(n1070), .A2(\completionDataOut[1][54] ), .B1(n1084), 
        .B2(\completionDataOut[3][54] ), .ZN(n1787) );
  AOI22D1 U2085 ( .A1(n1045), .A2(\completionDataOut[0][54] ), .B1(n1058), 
        .B2(\completionDataOut[2][54] ), .ZN(n1786) );
  AOI22D1 U2086 ( .A1(n1120), .A2(\completionDataOut[5][53] ), .B1(n1134), 
        .B2(\completionDataOut[7][53] ), .ZN(n1785) );
  CKBD1 U2087 ( .I(n1142), .Z(n1134) );
  AOI22D1 U2088 ( .A1(n1096), .A2(\completionDataOut[4][53] ), .B1(n1109), 
        .B2(\completionDataOut[6][53] ), .ZN(n1784) );
  CKBD1 U2089 ( .I(n1117), .Z(n1109) );
  AOI22D1 U2090 ( .A1(n1070), .A2(\completionDataOut[1][53] ), .B1(n1084), 
        .B2(\completionDataOut[3][53] ), .ZN(n1783) );
  CKBD1 U2091 ( .I(n1092), .Z(n1084) );
  CKBD1 U2092 ( .I(n1082), .Z(n1070) );
  AOI22D1 U2093 ( .A1(n1045), .A2(\completionDataOut[0][53] ), .B1(n1058), 
        .B2(\completionDataOut[2][53] ), .ZN(n1782) );
  CKBD1 U2094 ( .I(n1066), .Z(n1058) );
  CKBD1 U2095 ( .I(n492), .Z(n1045) );
  AOI22D1 U2096 ( .A1(n1046), .A2(\completionDataOut[0][52] ), .B1(n1067), 
        .B2(\completionDataOut[2][52] ), .ZN(n1780) );
  AOI22D1 U2097 ( .A1(n1046), .A2(\completionDataOut[0][51] ), .B1(n1066), 
        .B2(\completionDataOut[2][51] ), .ZN(n1779) );
  AOI22D1 U2098 ( .A1(n1121), .A2(\completionDataOut[5][50] ), .B1(n1142), 
        .B2(\completionDataOut[7][50] ), .ZN(n1778) );
  AOI22D1 U2099 ( .A1(n1097), .A2(\completionDataOut[4][50] ), .B1(n1117), 
        .B2(\completionDataOut[6][50] ), .ZN(n1777) );
  AOI22D1 U2100 ( .A1(n1071), .A2(\completionDataOut[1][50] ), .B1(n1092), 
        .B2(\completionDataOut[3][50] ), .ZN(n1776) );
  AOI22D1 U2101 ( .A1(n1046), .A2(\completionDataOut[0][50] ), .B1(n1066), 
        .B2(\completionDataOut[2][50] ), .ZN(n1775) );
  AOI22D1 U2102 ( .A1(n1121), .A2(\completionDataOut[5][49] ), .B1(n1142), 
        .B2(\completionDataOut[7][49] ), .ZN(n1774) );
  AOI22D1 U2103 ( .A1(n1097), .A2(\completionDataOut[4][49] ), .B1(n1117), 
        .B2(\completionDataOut[6][49] ), .ZN(n1773) );
  AOI22D1 U2104 ( .A1(n1071), .A2(\completionDataOut[1][49] ), .B1(n1092), 
        .B2(\completionDataOut[3][49] ), .ZN(n1772) );
  AOI22D1 U2105 ( .A1(n1046), .A2(\completionDataOut[0][49] ), .B1(n1066), 
        .B2(\completionDataOut[2][49] ), .ZN(n1771) );
  AOI22D1 U2106 ( .A1(n1121), .A2(\completionDataOut[5][48] ), .B1(n1143), 
        .B2(\completionDataOut[7][48] ), .ZN(n1770) );
  AOI22D1 U2107 ( .A1(n1097), .A2(\completionDataOut[4][48] ), .B1(n1118), 
        .B2(\completionDataOut[6][48] ), .ZN(n1769) );
  AOI22D1 U2108 ( .A1(n1071), .A2(\completionDataOut[1][48] ), .B1(n1093), 
        .B2(\completionDataOut[3][48] ), .ZN(n1768) );
  AOI22D1 U2109 ( .A1(n1046), .A2(\completionDataOut[0][48] ), .B1(n1067), 
        .B2(\completionDataOut[2][48] ), .ZN(n1767) );
  AOI22D1 U2110 ( .A1(n1121), .A2(\completionDataOut[5][47] ), .B1(n1143), 
        .B2(\completionDataOut[7][47] ), .ZN(n1766) );
  AOI22D1 U2111 ( .A1(n1097), .A2(\completionDataOut[4][47] ), .B1(n1118), 
        .B2(\completionDataOut[6][47] ), .ZN(n1765) );
  AOI22D1 U2112 ( .A1(n1071), .A2(\completionDataOut[1][47] ), .B1(n1093), 
        .B2(\completionDataOut[3][47] ), .ZN(n1764) );
  CKBD1 U2113 ( .I(n1080), .Z(n1071) );
  AOI22D1 U2114 ( .A1(n1046), .A2(\completionDataOut[0][47] ), .B1(n1067), 
        .B2(\completionDataOut[2][47] ), .ZN(n1763) );
  CKBD1 U2115 ( .I(n1055), .Z(n1046) );
  AOI22D1 U2116 ( .A1(n1072), .A2(\completionDataOut[1][46] ), .B1(n1085), 
        .B2(\completionDataOut[3][46] ), .ZN(n1760) );
  AOI22D1 U2117 ( .A1(n1047), .A2(\completionDataOut[0][46] ), .B1(n1059), 
        .B2(\completionDataOut[2][46] ), .ZN(n1759) );
  AOI22D1 U2118 ( .A1(n1072), .A2(\completionDataOut[1][45] ), .B1(n1085), 
        .B2(\completionDataOut[3][45] ), .ZN(n1757) );
  AOI22D1 U2119 ( .A1(n1047), .A2(\completionDataOut[0][45] ), .B1(n1059), 
        .B2(\completionDataOut[2][45] ), .ZN(n1756) );
  AOI22D1 U2120 ( .A1(n1098), .A2(\completionDataOut[4][44] ), .B1(n1110), 
        .B2(\completionDataOut[6][44] ), .ZN(n1755) );
  AOI22D1 U2121 ( .A1(n1122), .A2(\completionDataOut[5][43] ), .B1(n1135), 
        .B2(\completionDataOut[7][43] ), .ZN(n1754) );
  AOI22D1 U2122 ( .A1(n1098), .A2(\completionDataOut[4][43] ), .B1(n1110), 
        .B2(\completionDataOut[6][43] ), .ZN(n1753) );
  AOI22D1 U2123 ( .A1(n1072), .A2(\completionDataOut[1][43] ), .B1(n1085), 
        .B2(\completionDataOut[3][43] ), .ZN(n1752) );
  AOI22D1 U2124 ( .A1(n1047), .A2(\completionDataOut[0][43] ), .B1(n1059), 
        .B2(\completionDataOut[2][43] ), .ZN(n1751) );
  AOI22D1 U2125 ( .A1(n1122), .A2(\completionDataOut[5][42] ), .B1(n1135), 
        .B2(\completionDataOut[7][42] ), .ZN(n1750) );
  AOI22D1 U2126 ( .A1(n1072), .A2(\completionDataOut[1][42] ), .B1(n1085), 
        .B2(\completionDataOut[3][42] ), .ZN(n1748) );
  AOI22D1 U2127 ( .A1(n1047), .A2(\completionDataOut[0][42] ), .B1(n1059), 
        .B2(\completionDataOut[2][42] ), .ZN(n1747) );
  AOI22D1 U2128 ( .A1(n1122), .A2(\completionDataOut[5][41] ), .B1(n1135), 
        .B2(\completionDataOut[7][41] ), .ZN(n1746) );
  CKBD1 U2129 ( .I(n1141), .Z(n1135) );
  AOI22D1 U2130 ( .A1(n1098), .A2(\completionDataOut[4][41] ), .B1(n1110), 
        .B2(\completionDataOut[6][41] ), .ZN(n1745) );
  CKBD1 U2131 ( .I(n1116), .Z(n1110) );
  AOI22D1 U2132 ( .A1(n1072), .A2(\completionDataOut[1][41] ), .B1(n1085), 
        .B2(\completionDataOut[3][41] ), .ZN(n1744) );
  CKBD1 U2133 ( .I(n1091), .Z(n1085) );
  CKBD1 U2134 ( .I(n1080), .Z(n1072) );
  AOI22D1 U2135 ( .A1(n1047), .A2(\completionDataOut[0][41] ), .B1(n1059), 
        .B2(\completionDataOut[2][41] ), .ZN(n1743) );
  CKBD1 U2136 ( .I(n1065), .Z(n1059) );
  CKBD1 U2137 ( .I(n1055), .Z(n1047) );
  AOI22D1 U2138 ( .A1(n1073), .A2(\completionDataOut[1][40] ), .B1(n1093), 
        .B2(\completionDataOut[3][40] ), .ZN(n1740) );
  AOI22D1 U2139 ( .A1(n1048), .A2(\completionDataOut[0][40] ), .B1(n1067), 
        .B2(\completionDataOut[2][40] ), .ZN(n1739) );
  AOI22D1 U2140 ( .A1(n1073), .A2(\completionDataOut[1][39] ), .B1(n1091), 
        .B2(\completionDataOut[3][39] ), .ZN(n1738) );
  AOI22D1 U2141 ( .A1(n1048), .A2(\completionDataOut[0][39] ), .B1(n1065), 
        .B2(\completionDataOut[2][39] ), .ZN(n1737) );
  AOI22D1 U2142 ( .A1(n1048), .A2(\completionDataOut[0][38] ), .B1(n1065), 
        .B2(\completionDataOut[2][38] ), .ZN(n1736) );
  AOI22D1 U2143 ( .A1(n1123), .A2(\completionDataOut[5][37] ), .B1(n1141), 
        .B2(\completionDataOut[7][37] ), .ZN(n1735) );
  AOI22D1 U2144 ( .A1(n1099), .A2(\completionDataOut[4][37] ), .B1(n1116), 
        .B2(\completionDataOut[6][37] ), .ZN(n1734) );
  AOI22D1 U2145 ( .A1(n1073), .A2(\completionDataOut[1][37] ), .B1(n1091), 
        .B2(\completionDataOut[3][37] ), .ZN(n1733) );
  AOI22D1 U2146 ( .A1(n1048), .A2(\completionDataOut[0][37] ), .B1(n1065), 
        .B2(\completionDataOut[2][37] ), .ZN(n1732) );
  AOI22D1 U2147 ( .A1(n1123), .A2(\completionDataOut[5][36] ), .B1(n1141), 
        .B2(\completionDataOut[7][36] ), .ZN(n1731) );
  AOI22D1 U2148 ( .A1(n1099), .A2(\completionDataOut[4][36] ), .B1(n1116), 
        .B2(\completionDataOut[6][36] ), .ZN(n1730) );
  AOI22D1 U2149 ( .A1(n1073), .A2(\completionDataOut[1][36] ), .B1(n1091), 
        .B2(\completionDataOut[3][36] ), .ZN(n1729) );
  AOI22D1 U2150 ( .A1(n1048), .A2(\completionDataOut[0][36] ), .B1(n1065), 
        .B2(\completionDataOut[2][36] ), .ZN(n1728) );
  AOI22D1 U2151 ( .A1(n1123), .A2(\completionDataOut[5][35] ), .B1(n1141), 
        .B2(\completionDataOut[7][35] ), .ZN(n1727) );
  AOI22D1 U2152 ( .A1(n1099), .A2(\completionDataOut[4][35] ), .B1(n1116), 
        .B2(\completionDataOut[6][35] ), .ZN(n1726) );
  AOI22D1 U2153 ( .A1(n1073), .A2(\completionDataOut[1][35] ), .B1(n1091), 
        .B2(\completionDataOut[3][35] ), .ZN(n1725) );
  CKBD1 U2154 ( .I(n1082), .Z(n1073) );
  AOI22D1 U2155 ( .A1(n1048), .A2(\completionDataOut[0][35] ), .B1(n1065), 
        .B2(\completionDataOut[2][35] ), .ZN(n1724) );
  CKBD1 U2156 ( .I(n1067), .Z(n1065) );
  CKBD1 U2157 ( .I(n492), .Z(n1048) );
  AOI22D1 U2158 ( .A1(n1074), .A2(\completionDataOut[1][34] ), .B1(n1086), 
        .B2(\completionDataOut[3][34] ), .ZN(n1721) );
  AOI22D1 U2159 ( .A1(n1049), .A2(\completionDataOut[0][34] ), .B1(n1060), 
        .B2(\completionDataOut[2][34] ), .ZN(n1720) );
  AOI22D1 U2160 ( .A1(n1074), .A2(\completionDataOut[1][33] ), .B1(n1086), 
        .B2(\completionDataOut[3][33] ), .ZN(n1717) );
  AOI22D1 U2161 ( .A1(n1049), .A2(\completionDataOut[0][33] ), .B1(n1060), 
        .B2(\completionDataOut[2][33] ), .ZN(n1716) );
  AOI22D1 U2162 ( .A1(n1074), .A2(\completionDataOut[1][32] ), .B1(n1086), 
        .B2(\completionDataOut[3][32] ), .ZN(n1713) );
  AOI22D1 U2163 ( .A1(n1049), .A2(\completionDataOut[0][32] ), .B1(n1060), 
        .B2(\completionDataOut[2][32] ), .ZN(n1712) );
  AOI22D1 U2164 ( .A1(n1124), .A2(\completionDataOut[5][31] ), .B1(n1136), 
        .B2(\completionDataOut[7][31] ), .ZN(n1711) );
  AOI22D1 U2165 ( .A1(n1100), .A2(\completionDataOut[4][31] ), .B1(n1111), 
        .B2(\completionDataOut[6][31] ), .ZN(n1710) );
  AOI22D1 U2166 ( .A1(n1074), .A2(\completionDataOut[1][31] ), .B1(n1086), 
        .B2(\completionDataOut[3][31] ), .ZN(n1709) );
  AOI22D1 U2167 ( .A1(n1049), .A2(\completionDataOut[0][31] ), .B1(n1060), 
        .B2(\completionDataOut[2][31] ), .ZN(n1708) );
  AOI22D1 U2168 ( .A1(n1074), .A2(\completionDataOut[1][30] ), .B1(n1086), 
        .B2(\completionDataOut[3][30] ), .ZN(n1707) );
  AOI22D1 U2169 ( .A1(n1049), .A2(\completionDataOut[0][30] ), .B1(n1060), 
        .B2(\completionDataOut[2][30] ), .ZN(n1706) );
  AOI22D1 U2170 ( .A1(n1124), .A2(\completionDataOut[5][29] ), .B1(n1136), 
        .B2(\completionDataOut[7][29] ), .ZN(n1705) );
  CKBD1 U2171 ( .I(n1144), .Z(n1136) );
  CKBD1 U2172 ( .I(n1129), .Z(n1124) );
  AOI22D1 U2173 ( .A1(n1100), .A2(\completionDataOut[4][29] ), .B1(n1111), 
        .B2(\completionDataOut[6][29] ), .ZN(n1704) );
  CKBD1 U2174 ( .I(n1119), .Z(n1111) );
  CKBD1 U2175 ( .I(n1105), .Z(n1100) );
  AOI22D1 U2176 ( .A1(n1074), .A2(\completionDataOut[1][29] ), .B1(n1086), 
        .B2(\completionDataOut[3][29] ), .ZN(n1703) );
  CKBD1 U2177 ( .I(n1094), .Z(n1086) );
  CKBD1 U2178 ( .I(n1079), .Z(n1074) );
  AOI22D1 U2179 ( .A1(n1049), .A2(\completionDataOut[0][29] ), .B1(n1060), 
        .B2(\completionDataOut[2][29] ), .ZN(n1702) );
  CKBD1 U2180 ( .I(n1068), .Z(n1060) );
  CKBD1 U2181 ( .I(n1054), .Z(n1049) );
  AOI22D1 U2182 ( .A1(n1081), .A2(\completionDataOut[1][28] ), .B1(n1087), 
        .B2(\completionDataOut[3][28] ), .ZN(n1701) );
  AOI22D1 U2183 ( .A1(n1056), .A2(\completionDataOut[0][28] ), .B1(n1061), 
        .B2(\completionDataOut[2][28] ), .ZN(n1700) );
  AOI22D1 U2184 ( .A1(n1079), .A2(\completionDataOut[1][27] ), .B1(n1087), 
        .B2(\completionDataOut[3][27] ), .ZN(n1697) );
  AOI22D1 U2185 ( .A1(n1054), .A2(\completionDataOut[0][27] ), .B1(n1061), 
        .B2(\completionDataOut[2][27] ), .ZN(n1696) );
  AOI22D1 U2186 ( .A1(n1079), .A2(\completionDataOut[1][26] ), .B1(n1087), 
        .B2(\completionDataOut[3][26] ), .ZN(n1693) );
  AOI22D1 U2187 ( .A1(n1054), .A2(\completionDataOut[0][26] ), .B1(n1061), 
        .B2(\completionDataOut[2][26] ), .ZN(n1692) );
  AOI22D1 U2188 ( .A1(n1054), .A2(\completionDataOut[0][25] ), .B1(n1061), 
        .B2(\completionDataOut[2][25] ), .ZN(n1691) );
  AOI22D1 U2189 ( .A1(n1129), .A2(\completionDataOut[5][24] ), .B1(n1137), 
        .B2(\completionDataOut[7][24] ), .ZN(n1690) );
  AOI22D1 U2190 ( .A1(n1105), .A2(\completionDataOut[4][24] ), .B1(n1112), 
        .B2(\completionDataOut[6][24] ), .ZN(n1689) );
  AOI22D1 U2191 ( .A1(n1079), .A2(\completionDataOut[1][24] ), .B1(n1087), 
        .B2(\completionDataOut[3][24] ), .ZN(n1688) );
  AOI22D1 U2192 ( .A1(n1054), .A2(\completionDataOut[0][24] ), .B1(n1061), 
        .B2(\completionDataOut[2][24] ), .ZN(n1687) );
  AOI22D1 U2193 ( .A1(n1129), .A2(\completionDataOut[5][23] ), .B1(n1137), 
        .B2(\completionDataOut[7][23] ), .ZN(n1686) );
  CKBD1 U2194 ( .I(n1131), .Z(n1129) );
  AOI22D1 U2195 ( .A1(n1105), .A2(\completionDataOut[4][23] ), .B1(n1112), 
        .B2(\completionDataOut[6][23] ), .ZN(n1685) );
  CKBD1 U2196 ( .I(n1107), .Z(n1105) );
  AOI22D1 U2197 ( .A1(n1079), .A2(\completionDataOut[1][23] ), .B1(n1087), 
        .B2(\completionDataOut[3][23] ), .ZN(n1684) );
  CKBD1 U2198 ( .I(n1081), .Z(n1079) );
  AOI22D1 U2199 ( .A1(n1054), .A2(\completionDataOut[0][23] ), .B1(n1061), 
        .B2(\completionDataOut[2][23] ), .ZN(n1683) );
  CKBD1 U2200 ( .I(n1069), .Z(n1061) );
  CKBD1 U2201 ( .I(n1056), .Z(n1054) );
  AOI22D1 U2202 ( .A1(n1075), .A2(\completionDataOut[1][22] ), .B1(n1088), 
        .B2(\completionDataOut[3][22] ), .ZN(n1680) );
  AOI22D1 U2203 ( .A1(n1050), .A2(\completionDataOut[0][22] ), .B1(n1062), 
        .B2(\completionDataOut[2][22] ), .ZN(n1679) );
  AOI22D1 U2204 ( .A1(n1075), .A2(\completionDataOut[1][21] ), .B1(n1088), 
        .B2(\completionDataOut[3][21] ), .ZN(n1676) );
  AOI22D1 U2205 ( .A1(n1050), .A2(\completionDataOut[0][21] ), .B1(n1062), 
        .B2(\completionDataOut[2][21] ), .ZN(n1675) );
  AOI22D1 U2206 ( .A1(n1075), .A2(\completionDataOut[1][20] ), .B1(n1088), 
        .B2(\completionDataOut[3][20] ), .ZN(n1672) );
  AOI22D1 U2207 ( .A1(n1050), .A2(\completionDataOut[0][20] ), .B1(n1062), 
        .B2(\completionDataOut[2][20] ), .ZN(n1671) );
  AOI22D1 U2208 ( .A1(n1125), .A2(\completionDataOut[5][19] ), .B1(n1138), 
        .B2(\completionDataOut[7][19] ), .ZN(n1670) );
  AOI22D1 U2209 ( .A1(n1101), .A2(\completionDataOut[4][19] ), .B1(n1113), 
        .B2(\completionDataOut[6][19] ), .ZN(n1669) );
  AOI22D1 U2210 ( .A1(n1075), .A2(\completionDataOut[1][19] ), .B1(n1088), 
        .B2(\completionDataOut[3][19] ), .ZN(n1668) );
  AOI22D1 U2211 ( .A1(n1050), .A2(\completionDataOut[0][19] ), .B1(n1062), 
        .B2(\completionDataOut[2][19] ), .ZN(n1667) );
  AOI22D1 U2212 ( .A1(n1101), .A2(\completionDataOut[4][18] ), .B1(n1113), 
        .B2(\completionDataOut[6][18] ), .ZN(n1666) );
  AOI22D1 U2213 ( .A1(n1050), .A2(\completionDataOut[0][18] ), .B1(n1062), 
        .B2(\completionDataOut[2][18] ), .ZN(n1665) );
  AOI22D1 U2214 ( .A1(n1125), .A2(\completionDataOut[5][17] ), .B1(n1138), 
        .B2(\completionDataOut[7][17] ), .ZN(n1664) );
  CKBD1 U2215 ( .I(n1140), .Z(n1138) );
  CKBD1 U2216 ( .I(n1128), .Z(n1125) );
  AOI22D1 U2217 ( .A1(n1101), .A2(\completionDataOut[4][17] ), .B1(n1113), 
        .B2(\completionDataOut[6][17] ), .ZN(n1663) );
  CKBD1 U2218 ( .I(n1115), .Z(n1113) );
  CKBD1 U2219 ( .I(n1104), .Z(n1101) );
  AOI22D1 U2220 ( .A1(n1075), .A2(\completionDataOut[1][17] ), .B1(n1088), 
        .B2(\completionDataOut[3][17] ), .ZN(n1662) );
  CKBD1 U2221 ( .I(n1090), .Z(n1088) );
  AOI22D1 U2222 ( .A1(n1050), .A2(\completionDataOut[0][17] ), .B1(n1062), 
        .B2(\completionDataOut[2][17] ), .ZN(n1661) );
  CKBD1 U2223 ( .I(n1064), .Z(n1062) );
  CKBD1 U2224 ( .I(n1053), .Z(n1050) );
  AOI22D1 U2225 ( .A1(n1078), .A2(\completionDataOut[1][16] ), .B1(n1095), 
        .B2(\completionDataOut[3][16] ), .ZN(n1658) );
  AOI22D1 U2226 ( .A1(n1053), .A2(\completionDataOut[0][16] ), .B1(n1069), 
        .B2(\completionDataOut[2][16] ), .ZN(n1657) );
  AOI22D1 U2227 ( .A1(n1131), .A2(\completionDataOut[5][15] ), .B1(n1145), 
        .B2(\completionDataOut[7][15] ), .ZN(n1656) );
  AOI22D1 U2228 ( .A1(n1107), .A2(\completionDataOut[4][15] ), .B1(n1601), 
        .B2(\completionDataOut[6][15] ), .ZN(n1655) );
  AOI22D1 U2229 ( .A1(n1081), .A2(\completionDataOut[1][15] ), .B1(n1095), 
        .B2(\completionDataOut[3][15] ), .ZN(n1654) );
  AOI22D1 U2230 ( .A1(n1056), .A2(\completionDataOut[0][15] ), .B1(n1069), 
        .B2(\completionDataOut[2][15] ), .ZN(n1653) );
  AOI22D1 U2231 ( .A1(n1078), .A2(\completionDataOut[1][14] ), .B1(n1094), 
        .B2(\completionDataOut[3][14] ), .ZN(n1650) );
  AOI22D1 U2232 ( .A1(n1053), .A2(\completionDataOut[0][14] ), .B1(n1068), 
        .B2(\completionDataOut[2][14] ), .ZN(n1649) );
  AOI22D1 U2233 ( .A1(n1053), .A2(\completionDataOut[0][13] ), .B1(n1068), 
        .B2(\completionDataOut[2][13] ), .ZN(n1648) );
  AOI22D1 U2234 ( .A1(n1128), .A2(\completionDataOut[5][12] ), .B1(n1144), 
        .B2(\completionDataOut[7][12] ), .ZN(n1647) );
  AOI22D1 U2235 ( .A1(n1104), .A2(\completionDataOut[4][12] ), .B1(n1119), 
        .B2(\completionDataOut[6][12] ), .ZN(n1646) );
  AOI22D1 U2236 ( .A1(n1078), .A2(\completionDataOut[1][12] ), .B1(n1094), 
        .B2(\completionDataOut[3][12] ), .ZN(n1645) );
  AOI22D1 U2237 ( .A1(n1053), .A2(\completionDataOut[0][12] ), .B1(n1068), 
        .B2(\completionDataOut[2][12] ), .ZN(n1644) );
  AOI22D1 U2238 ( .A1(n1128), .A2(\completionDataOut[5][11] ), .B1(n1144), 
        .B2(\completionDataOut[7][11] ), .ZN(n1643) );
  CKBD1 U2239 ( .I(n1131), .Z(n1128) );
  AOI22D1 U2240 ( .A1(n1104), .A2(\completionDataOut[4][11] ), .B1(n1119), 
        .B2(\completionDataOut[6][11] ), .ZN(n1642) );
  CKBD1 U2241 ( .I(n1107), .Z(n1104) );
  AOI22D1 U2242 ( .A1(n1078), .A2(\completionDataOut[1][11] ), .B1(n1094), 
        .B2(\completionDataOut[3][11] ), .ZN(n1641) );
  CKBD1 U2243 ( .I(n1081), .Z(n1078) );
  AOI22D1 U2244 ( .A1(n1053), .A2(\completionDataOut[0][11] ), .B1(n1068), 
        .B2(\completionDataOut[2][11] ), .ZN(n1640) );
  CKBD1 U2245 ( .I(n1056), .Z(n1053) );
  AOI22D1 U2246 ( .A1(n1077), .A2(\completionDataOut[1][10] ), .B1(n1089), 
        .B2(\completionDataOut[3][10] ), .ZN(n1637) );
  AOI22D1 U2247 ( .A1(n1052), .A2(\completionDataOut[0][10] ), .B1(n1063), 
        .B2(\completionDataOut[2][10] ), .ZN(n1636) );
  AOI22D1 U2248 ( .A1(n1077), .A2(\completionDataOut[1][9] ), .B1(n1089), .B2(
        \completionDataOut[3][9] ), .ZN(n1635) );
  AOI22D1 U2249 ( .A1(n1052), .A2(\completionDataOut[0][9] ), .B1(n1063), .B2(
        \completionDataOut[2][9] ), .ZN(n1634) );
  AOI22D1 U2250 ( .A1(n1127), .A2(\completionDataOut[5][8] ), .B1(n1139), .B2(
        \completionDataOut[7][8] ), .ZN(n1633) );
  AOI22D1 U2251 ( .A1(n1103), .A2(\completionDataOut[4][8] ), .B1(n1114), .B2(
        \completionDataOut[6][8] ), .ZN(n1632) );
  AOI22D1 U2252 ( .A1(n1077), .A2(\completionDataOut[1][8] ), .B1(n1089), .B2(
        \completionDataOut[3][8] ), .ZN(n1631) );
  AOI22D1 U2253 ( .A1(n1052), .A2(\completionDataOut[0][8] ), .B1(n1063), .B2(
        \completionDataOut[2][8] ), .ZN(n1630) );
  CKBD1 U2254 ( .I(n1142), .Z(n1133) );
  CKBD1 U2255 ( .I(n1117), .Z(n1108) );
  AOI22D1 U2256 ( .A1(n1080), .A2(\completionDataOut[1][62] ), .B1(n1083), 
        .B2(\completionDataOut[3][62] ), .ZN(n1813) );
  CKBD1 U2257 ( .I(n1092), .Z(n1083) );
  CKBD1 U2258 ( .I(n1066), .Z(n1057) );
  CKBD1 U2259 ( .I(n1067), .Z(n1066) );
  AOI22D1 U2260 ( .A1(n1127), .A2(\completionDataOut[5][7] ), .B1(n1139), .B2(
        \completionDataOut[7][7] ), .ZN(n1629) );
  AOI22D1 U2261 ( .A1(n1103), .A2(\completionDataOut[4][7] ), .B1(n1114), .B2(
        \completionDataOut[6][7] ), .ZN(n1628) );
  AOI22D1 U2262 ( .A1(n1077), .A2(\completionDataOut[1][7] ), .B1(n1089), .B2(
        \completionDataOut[3][7] ), .ZN(n1627) );
  AOI22D1 U2263 ( .A1(n1052), .A2(\completionDataOut[0][7] ), .B1(n1063), .B2(
        \completionDataOut[2][7] ), .ZN(n1626) );
  AOI22D1 U2264 ( .A1(n1127), .A2(\completionDataOut[5][6] ), .B1(n1139), .B2(
        \completionDataOut[7][6] ), .ZN(n1625) );
  AOI22D1 U2265 ( .A1(n1077), .A2(\completionDataOut[1][6] ), .B1(n1089), .B2(
        \completionDataOut[3][6] ), .ZN(n1623) );
  AOI22D1 U2266 ( .A1(n1052), .A2(\completionDataOut[0][6] ), .B1(n1063), .B2(
        \completionDataOut[2][6] ), .ZN(n1622) );
  AOI22D1 U2267 ( .A1(n1051), .A2(\completionDataOut[0][5] ), .B1(n1063), .B2(
        \completionDataOut[2][5] ), .ZN(n1621) );
  CKBD1 U2268 ( .I(n1069), .Z(n1063) );
  AOI22D1 U2269 ( .A1(n1051), .A2(\completionDataOut[0][4] ), .B1(n1064), .B2(
        \completionDataOut[2][4] ), .ZN(n1620) );
  AOI22D1 U2270 ( .A1(n1126), .A2(\completionDataOut[5][3] ), .B1(n1140), .B2(
        \completionDataOut[7][3] ), .ZN(n1619) );
  AOI22D1 U2271 ( .A1(n1102), .A2(\completionDataOut[4][3] ), .B1(n1115), .B2(
        \completionDataOut[6][3] ), .ZN(n1618) );
  AOI22D1 U2272 ( .A1(n1076), .A2(\completionDataOut[1][3] ), .B1(n1090), .B2(
        \completionDataOut[3][3] ), .ZN(n1617) );
  AOI22D1 U2273 ( .A1(n1051), .A2(\completionDataOut[0][3] ), .B1(n1064), .B2(
        \completionDataOut[2][3] ), .ZN(n1616) );
  AOI22D1 U2274 ( .A1(n1126), .A2(\completionDataOut[5][2] ), .B1(n1140), .B2(
        \completionDataOut[7][2] ), .ZN(n1615) );
  AOI22D1 U2275 ( .A1(n1102), .A2(\completionDataOut[4][2] ), .B1(n1115), .B2(
        \completionDataOut[6][2] ), .ZN(n1614) );
  AOI22D1 U2276 ( .A1(n1076), .A2(\completionDataOut[1][2] ), .B1(n1090), .B2(
        \completionDataOut[3][2] ), .ZN(n1613) );
  AOI22D1 U2277 ( .A1(n1051), .A2(\completionDataOut[0][2] ), .B1(n1064), .B2(
        \completionDataOut[2][2] ), .ZN(n1612) );
  AOI22D1 U2278 ( .A1(n1126), .A2(\completionDataOut[5][1] ), .B1(n1140), .B2(
        \completionDataOut[7][1] ), .ZN(n1611) );
  AOI22D1 U2279 ( .A1(n1102), .A2(\completionDataOut[4][1] ), .B1(n1115), .B2(
        \completionDataOut[6][1] ), .ZN(n1610) );
  AOI22D1 U2280 ( .A1(n1076), .A2(\completionDataOut[1][1] ), .B1(n1090), .B2(
        \completionDataOut[3][1] ), .ZN(n1609) );
  AOI22D1 U2281 ( .A1(n1051), .A2(\completionDataOut[0][1] ), .B1(n1064), .B2(
        \completionDataOut[2][1] ), .ZN(n1608) );
  AOI22D1 U2282 ( .A1(n1126), .A2(\completionDataOut[5][0] ), .B1(n1140), .B2(
        \completionDataOut[7][0] ), .ZN(n1607) );
  CKBD1 U2283 ( .I(n1131), .Z(n1127) );
  AOI22D1 U2284 ( .A1(n1102), .A2(\completionDataOut[4][0] ), .B1(n1115), .B2(
        \completionDataOut[6][0] ), .ZN(n1606) );
  CKBD1 U2285 ( .I(n1107), .Z(n1103) );
  AOI22D1 U2286 ( .A1(n1076), .A2(\completionDataOut[1][0] ), .B1(n1090), .B2(
        \completionDataOut[3][0] ), .ZN(n1605) );
  NR2D1 U2287 ( .A1(decodeReadAddr1_i[2]), .A2(n1598), .ZN(n1599) );
  ND2D1 U2288 ( .A1(decodeReadAddr1_i[0]), .A2(decodeReadAddr1_i[1]), .ZN(
        n1598) );
  CKBD1 U2289 ( .I(n1081), .Z(n1077) );
  CKBD1 U2290 ( .I(n1082), .Z(n1081) );
  NR2D1 U2291 ( .A1(decodeReadAddr1_i[2]), .A2(n1596), .ZN(n1597) );
  INVD1 U2292 ( .I(decodeReadAddr1_i[1]), .ZN(n1823) );
  AOI22D1 U2293 ( .A1(n1051), .A2(\completionDataOut[0][0] ), .B1(n1064), .B2(
        \completionDataOut[2][0] ), .ZN(n1604) );
  CKBD1 U2294 ( .I(n1068), .Z(n1064) );
  NR2D1 U2295 ( .A1(decodeReadAddr1_i[2]), .A2(n1594), .ZN(n1595) );
  ND2D1 U2296 ( .A1(decodeReadAddr1_i[1]), .A2(n1822), .ZN(n1594) );
  INVD1 U2297 ( .I(decodeReadAddr1_i[0]), .ZN(n1822) );
  CKBD1 U2298 ( .I(n1052), .Z(n1051) );
  CKBD1 U2299 ( .I(n1056), .Z(n1052) );
  AOI22D1 U2300 ( .A1(n1183), .A2(\completionDataOut[1][64] ), .B1(n1184), 
        .B2(\completionDataOut[3][64] ), .ZN(n2055) );
  AOI22D1 U2301 ( .A1(n493), .A2(\completionDataOut[0][64] ), .B1(n1158), .B2(
        \completionDataOut[2][64] ), .ZN(n2054) );
  AOI22D1 U2302 ( .A1(n1183), .A2(\completionDataOut[1][63] ), .B1(n1184), 
        .B2(\completionDataOut[3][63] ), .ZN(n2051) );
  AOI22D1 U2303 ( .A1(n493), .A2(\completionDataOut[0][63] ), .B1(n1158), .B2(
        \completionDataOut[2][63] ), .ZN(n2050) );
  AOI22D1 U2304 ( .A1(n1232), .A2(\completionDataOut[5][62] ), .B1(n1234), 
        .B2(\completionDataOut[7][62] ), .ZN(n2049) );
  AOI22D1 U2305 ( .A1(n1207), .A2(\completionDataOut[4][62] ), .B1(n1209), 
        .B2(\completionDataOut[6][62] ), .ZN(n2048) );
  AOI22D1 U2306 ( .A1(n1181), .A2(\completionDataOut[1][62] ), .B1(n1184), 
        .B2(\completionDataOut[3][62] ), .ZN(n2047) );
  AOI22D1 U2307 ( .A1(n1156), .A2(\completionDataOut[0][62] ), .B1(n1158), 
        .B2(\completionDataOut[2][62] ), .ZN(n2046) );
  AOI22D1 U2308 ( .A1(n1232), .A2(\completionDataOut[5][61] ), .B1(n1234), 
        .B2(\completionDataOut[7][61] ), .ZN(n2045) );
  AOI22D1 U2309 ( .A1(n1207), .A2(\completionDataOut[4][61] ), .B1(n1209), 
        .B2(\completionDataOut[6][61] ), .ZN(n2044) );
  AOI22D1 U2310 ( .A1(n1181), .A2(\completionDataOut[1][61] ), .B1(n1184), 
        .B2(\completionDataOut[3][61] ), .ZN(n2043) );
  AOI22D1 U2311 ( .A1(n1156), .A2(\completionDataOut[0][61] ), .B1(n1158), 
        .B2(\completionDataOut[2][61] ), .ZN(n2042) );
  AOI22D1 U2312 ( .A1(n1207), .A2(\completionDataOut[4][60] ), .B1(n1209), 
        .B2(\completionDataOut[6][60] ), .ZN(n2041) );
  CKBD1 U2313 ( .I(n1243), .Z(n1234) );
  CKBD1 U2314 ( .I(n1218), .Z(n1209) );
  AOI22D1 U2315 ( .A1(n1181), .A2(\completionDataOut[1][59] ), .B1(n1184), 
        .B2(\completionDataOut[3][59] ), .ZN(n2040) );
  CKBD1 U2316 ( .I(n1193), .Z(n1184) );
  AOI22D1 U2317 ( .A1(n1156), .A2(\completionDataOut[0][59] ), .B1(n1158), 
        .B2(\completionDataOut[2][59] ), .ZN(n2039) );
  CKBD1 U2318 ( .I(n1167), .Z(n1158) );
  AOI22D1 U2319 ( .A1(n1171), .A2(\completionDataOut[1][58] ), .B1(n1185), 
        .B2(\completionDataOut[3][58] ), .ZN(n2036) );
  AOI22D1 U2320 ( .A1(n1146), .A2(\completionDataOut[0][58] ), .B1(n1159), 
        .B2(\completionDataOut[2][58] ), .ZN(n2035) );
  AOI22D1 U2321 ( .A1(n1224), .A2(\completionDataOut[5][43] ), .B1(n1236), 
        .B2(\completionDataOut[7][43] ), .ZN(n1985) );
  AOI22D1 U2322 ( .A1(n1199), .A2(\completionDataOut[4][43] ), .B1(n1211), 
        .B2(\completionDataOut[6][43] ), .ZN(n1984) );
  AOI22D1 U2323 ( .A1(n1173), .A2(\completionDataOut[1][43] ), .B1(n1186), 
        .B2(\completionDataOut[3][43] ), .ZN(n1983) );
  AOI22D1 U2324 ( .A1(n1148), .A2(\completionDataOut[0][43] ), .B1(n1160), 
        .B2(\completionDataOut[2][43] ), .ZN(n1982) );
  AOI22D1 U2325 ( .A1(n1197), .A2(\completionDataOut[4][57] ), .B1(n1210), 
        .B2(\completionDataOut[6][57] ), .ZN(n2033) );
  AOI22D1 U2326 ( .A1(n1171), .A2(\completionDataOut[1][57] ), .B1(n1185), 
        .B2(\completionDataOut[3][57] ), .ZN(n2032) );
  AOI22D1 U2327 ( .A1(n1146), .A2(\completionDataOut[0][57] ), .B1(n1159), 
        .B2(\completionDataOut[2][57] ), .ZN(n2031) );
  AOI22D1 U2328 ( .A1(n1197), .A2(\completionDataOut[4][56] ), .B1(n1210), 
        .B2(\completionDataOut[6][56] ), .ZN(n2029) );
  AOI22D1 U2329 ( .A1(n1171), .A2(\completionDataOut[1][56] ), .B1(n1185), 
        .B2(\completionDataOut[3][56] ), .ZN(n2028) );
  AOI22D1 U2330 ( .A1(n1146), .A2(\completionDataOut[0][56] ), .B1(n1159), 
        .B2(\completionDataOut[2][56] ), .ZN(n2027) );
  AOI22D1 U2331 ( .A1(n1222), .A2(\completionDataOut[5][55] ), .B1(n1235), 
        .B2(\completionDataOut[7][55] ), .ZN(n2026) );
  AOI22D1 U2332 ( .A1(n1197), .A2(\completionDataOut[4][55] ), .B1(n1210), 
        .B2(\completionDataOut[6][55] ), .ZN(n2025) );
  AOI22D1 U2333 ( .A1(n1171), .A2(\completionDataOut[1][55] ), .B1(n1185), 
        .B2(\completionDataOut[3][55] ), .ZN(n2024) );
  AOI22D1 U2334 ( .A1(n1146), .A2(\completionDataOut[0][55] ), .B1(n1159), 
        .B2(\completionDataOut[2][55] ), .ZN(n2023) );
  AOI22D1 U2335 ( .A1(n1222), .A2(\completionDataOut[5][54] ), .B1(n1235), 
        .B2(\completionDataOut[7][54] ), .ZN(n2022) );
  AOI22D1 U2336 ( .A1(n1197), .A2(\completionDataOut[4][54] ), .B1(n1210), 
        .B2(\completionDataOut[6][54] ), .ZN(n2021) );
  AOI22D1 U2337 ( .A1(n1171), .A2(\completionDataOut[1][54] ), .B1(n1185), 
        .B2(\completionDataOut[3][54] ), .ZN(n2020) );
  AOI22D1 U2338 ( .A1(n1146), .A2(\completionDataOut[0][54] ), .B1(n1159), 
        .B2(\completionDataOut[2][54] ), .ZN(n2019) );
  CKBD1 U2339 ( .I(n1243), .Z(n1235) );
  CKBD1 U2340 ( .I(n1218), .Z(n1210) );
  AOI22D1 U2341 ( .A1(n1171), .A2(\completionDataOut[1][53] ), .B1(n1185), 
        .B2(\completionDataOut[3][53] ), .ZN(n2018) );
  CKBD1 U2342 ( .I(n1193), .Z(n1185) );
  CKBD1 U2343 ( .I(n1183), .Z(n1171) );
  AOI22D1 U2344 ( .A1(n1146), .A2(\completionDataOut[0][53] ), .B1(n1159), 
        .B2(\completionDataOut[2][53] ), .ZN(n2017) );
  CKBD1 U2345 ( .I(n1167), .Z(n1159) );
  CKBD1 U2346 ( .I(n493), .Z(n1146) );
  AOI22D1 U2347 ( .A1(n1223), .A2(\completionDataOut[5][52] ), .B1(n1244), 
        .B2(\completionDataOut[7][52] ), .ZN(n2016) );
  AOI22D1 U2348 ( .A1(n1198), .A2(\completionDataOut[4][52] ), .B1(n1219), 
        .B2(\completionDataOut[6][52] ), .ZN(n2015) );
  AOI22D1 U2349 ( .A1(n1172), .A2(\completionDataOut[1][52] ), .B1(n1194), 
        .B2(\completionDataOut[3][52] ), .ZN(n2014) );
  AOI22D1 U2350 ( .A1(n1147), .A2(\completionDataOut[0][52] ), .B1(n1168), 
        .B2(\completionDataOut[2][52] ), .ZN(n2013) );
  AOI22D1 U2351 ( .A1(n1223), .A2(\completionDataOut[5][51] ), .B1(n1243), 
        .B2(\completionDataOut[7][51] ), .ZN(n2012) );
  AOI22D1 U2352 ( .A1(n1198), .A2(\completionDataOut[4][51] ), .B1(n1218), 
        .B2(\completionDataOut[6][51] ), .ZN(n2011) );
  AOI22D1 U2353 ( .A1(n1172), .A2(\completionDataOut[1][51] ), .B1(n1193), 
        .B2(\completionDataOut[3][51] ), .ZN(n2010) );
  AOI22D1 U2354 ( .A1(n1147), .A2(\completionDataOut[0][51] ), .B1(n1167), 
        .B2(\completionDataOut[2][51] ), .ZN(n2009) );
  AOI22D1 U2355 ( .A1(n1172), .A2(\completionDataOut[1][50] ), .B1(n1193), 
        .B2(\completionDataOut[3][50] ), .ZN(n2008) );
  AOI22D1 U2356 ( .A1(n1147), .A2(\completionDataOut[0][50] ), .B1(n1167), 
        .B2(\completionDataOut[2][50] ), .ZN(n2007) );
  AOI22D1 U2357 ( .A1(n1223), .A2(\completionDataOut[5][49] ), .B1(n1243), 
        .B2(\completionDataOut[7][49] ), .ZN(n2006) );
  CKBD1 U2358 ( .I(n1244), .Z(n1243) );
  AOI22D1 U2359 ( .A1(n1198), .A2(\completionDataOut[4][49] ), .B1(n1218), 
        .B2(\completionDataOut[6][49] ), .ZN(n2005) );
  CKBD1 U2360 ( .I(n1219), .Z(n1218) );
  AOI22D1 U2361 ( .A1(n1172), .A2(\completionDataOut[1][49] ), .B1(n1193), 
        .B2(\completionDataOut[3][49] ), .ZN(n2004) );
  CKBD1 U2362 ( .I(n1194), .Z(n1193) );
  AOI22D1 U2363 ( .A1(n1147), .A2(\completionDataOut[0][49] ), .B1(n1167), 
        .B2(\completionDataOut[2][49] ), .ZN(n2003) );
  CKBD1 U2364 ( .I(n1168), .Z(n1167) );
  AOI22D1 U2365 ( .A1(n1223), .A2(\completionDataOut[5][48] ), .B1(n1244), 
        .B2(\completionDataOut[7][48] ), .ZN(n2002) );
  AOI22D1 U2366 ( .A1(n1198), .A2(\completionDataOut[4][48] ), .B1(n1219), 
        .B2(\completionDataOut[6][48] ), .ZN(n2001) );
  AOI22D1 U2367 ( .A1(n1172), .A2(\completionDataOut[1][48] ), .B1(n1194), 
        .B2(\completionDataOut[3][48] ), .ZN(n2000) );
  AOI22D1 U2368 ( .A1(n1147), .A2(\completionDataOut[0][48] ), .B1(n1168), 
        .B2(\completionDataOut[2][48] ), .ZN(n1999) );
  CKBD1 U2369 ( .I(n1181), .Z(n1172) );
  AOI22D1 U2370 ( .A1(n1147), .A2(\completionDataOut[0][47] ), .B1(n1168), 
        .B2(\completionDataOut[2][47] ), .ZN(n1998) );
  CKBD1 U2371 ( .I(n1156), .Z(n1147) );
  AOI22D1 U2372 ( .A1(n1173), .A2(\completionDataOut[1][46] ), .B1(n1186), 
        .B2(\completionDataOut[3][46] ), .ZN(n1995) );
  AOI22D1 U2373 ( .A1(n1148), .A2(\completionDataOut[0][46] ), .B1(n1160), 
        .B2(\completionDataOut[2][46] ), .ZN(n1994) );
  AOI22D1 U2374 ( .A1(n1199), .A2(\completionDataOut[4][45] ), .B1(n1211), 
        .B2(\completionDataOut[6][45] ), .ZN(n1992) );
  AOI22D1 U2375 ( .A1(n1173), .A2(\completionDataOut[1][45] ), .B1(n1186), 
        .B2(\completionDataOut[3][45] ), .ZN(n1991) );
  AOI22D1 U2376 ( .A1(n1148), .A2(\completionDataOut[0][45] ), .B1(n1160), 
        .B2(\completionDataOut[2][45] ), .ZN(n1990) );
  AOI22D1 U2377 ( .A1(n1224), .A2(\completionDataOut[5][44] ), .B1(n1236), 
        .B2(\completionDataOut[7][44] ), .ZN(n1989) );
  AOI22D1 U2378 ( .A1(n1199), .A2(\completionDataOut[4][44] ), .B1(n1211), 
        .B2(\completionDataOut[6][44] ), .ZN(n1988) );
  AOI22D1 U2379 ( .A1(n1173), .A2(\completionDataOut[1][44] ), .B1(n1186), 
        .B2(\completionDataOut[3][44] ), .ZN(n1987) );
  AOI22D1 U2380 ( .A1(n1148), .A2(\completionDataOut[0][44] ), .B1(n1160), 
        .B2(\completionDataOut[2][44] ), .ZN(n1986) );
  AOI22D1 U2381 ( .A1(n1233), .A2(\completionDataOut[5][28] ), .B1(n1238), 
        .B2(\completionDataOut[7][28] ), .ZN(n1934) );
  AOI22D1 U2382 ( .A1(n1208), .A2(\completionDataOut[4][28] ), .B1(n1213), 
        .B2(\completionDataOut[6][28] ), .ZN(n1933) );
  AOI22D1 U2383 ( .A1(n1182), .A2(\completionDataOut[1][28] ), .B1(n1188), 
        .B2(\completionDataOut[3][28] ), .ZN(n1932) );
  AOI22D1 U2384 ( .A1(n1157), .A2(\completionDataOut[0][28] ), .B1(n1162), 
        .B2(\completionDataOut[2][28] ), .ZN(n1931) );
  AOI22D1 U2385 ( .A1(n1224), .A2(\completionDataOut[5][42] ), .B1(n1236), 
        .B2(\completionDataOut[7][42] ), .ZN(n1981) );
  AOI22D1 U2386 ( .A1(n1173), .A2(\completionDataOut[1][42] ), .B1(n1186), 
        .B2(\completionDataOut[3][42] ), .ZN(n1979) );
  AOI22D1 U2387 ( .A1(n1148), .A2(\completionDataOut[0][42] ), .B1(n1160), 
        .B2(\completionDataOut[2][42] ), .ZN(n1978) );
  CKBD1 U2388 ( .I(n1242), .Z(n1236) );
  CKBD1 U2389 ( .I(n1217), .Z(n1211) );
  AOI22D1 U2390 ( .A1(n1173), .A2(\completionDataOut[1][41] ), .B1(n1186), 
        .B2(\completionDataOut[3][41] ), .ZN(n1977) );
  CKBD1 U2391 ( .I(n1192), .Z(n1186) );
  CKBD1 U2392 ( .I(n1181), .Z(n1173) );
  AOI22D1 U2393 ( .A1(n1148), .A2(\completionDataOut[0][41] ), .B1(n1160), 
        .B2(\completionDataOut[2][41] ), .ZN(n1976) );
  CKBD1 U2394 ( .I(n1166), .Z(n1160) );
  CKBD1 U2395 ( .I(n1156), .Z(n1148) );
  AOI22D1 U2396 ( .A1(n1174), .A2(\completionDataOut[1][40] ), .B1(n1194), 
        .B2(\completionDataOut[3][40] ), .ZN(n1973) );
  AOI22D1 U2397 ( .A1(n1149), .A2(\completionDataOut[0][40] ), .B1(n1168), 
        .B2(\completionDataOut[2][40] ), .ZN(n1972) );
  AOI22D1 U2398 ( .A1(n1225), .A2(\completionDataOut[5][39] ), .B1(n1242), 
        .B2(\completionDataOut[7][39] ), .ZN(n1971) );
  AOI22D1 U2399 ( .A1(n1200), .A2(\completionDataOut[4][39] ), .B1(n1217), 
        .B2(\completionDataOut[6][39] ), .ZN(n1970) );
  AOI22D1 U2400 ( .A1(n1174), .A2(\completionDataOut[1][39] ), .B1(n1192), 
        .B2(\completionDataOut[3][39] ), .ZN(n1969) );
  AOI22D1 U2401 ( .A1(n1149), .A2(\completionDataOut[0][39] ), .B1(n1166), 
        .B2(\completionDataOut[2][39] ), .ZN(n1968) );
  AOI22D1 U2402 ( .A1(n1225), .A2(\completionDataOut[5][38] ), .B1(n1242), 
        .B2(\completionDataOut[7][38] ), .ZN(n1967) );
  AOI22D1 U2403 ( .A1(n1200), .A2(\completionDataOut[4][38] ), .B1(n1217), 
        .B2(\completionDataOut[6][38] ), .ZN(n1966) );
  AOI22D1 U2404 ( .A1(n1174), .A2(\completionDataOut[1][38] ), .B1(n1192), 
        .B2(\completionDataOut[3][38] ), .ZN(n1965) );
  AOI22D1 U2405 ( .A1(n1149), .A2(\completionDataOut[0][38] ), .B1(n1166), 
        .B2(\completionDataOut[2][38] ), .ZN(n1964) );
  AOI22D1 U2406 ( .A1(n1149), .A2(\completionDataOut[0][37] ), .B1(n1166), 
        .B2(\completionDataOut[2][37] ), .ZN(n1962) );
  AOI22D1 U2407 ( .A1(n1225), .A2(\completionDataOut[5][36] ), .B1(n1242), 
        .B2(\completionDataOut[7][36] ), .ZN(n1961) );
  AOI22D1 U2408 ( .A1(n1200), .A2(\completionDataOut[4][36] ), .B1(n1217), 
        .B2(\completionDataOut[6][36] ), .ZN(n1960) );
  AOI22D1 U2409 ( .A1(n1174), .A2(\completionDataOut[1][36] ), .B1(n1192), 
        .B2(\completionDataOut[3][36] ), .ZN(n1959) );
  AOI22D1 U2410 ( .A1(n1149), .A2(\completionDataOut[0][36] ), .B1(n1166), 
        .B2(\completionDataOut[2][36] ), .ZN(n1958) );
  CKBD1 U2411 ( .I(n1246), .Z(n1244) );
  CKBD1 U2412 ( .I(n1221), .Z(n1219) );
  AOI22D1 U2413 ( .A1(n1149), .A2(\completionDataOut[0][35] ), .B1(n1166), 
        .B2(\completionDataOut[2][35] ), .ZN(n1956) );
  CKBD1 U2414 ( .I(n1168), .Z(n1166) );
  CKBD1 U2415 ( .I(n493), .Z(n1149) );
  AOI22D1 U2416 ( .A1(n1175), .A2(\completionDataOut[1][34] ), .B1(n1187), 
        .B2(\completionDataOut[3][34] ), .ZN(n1953) );
  AOI22D1 U2417 ( .A1(n1150), .A2(\completionDataOut[0][34] ), .B1(n1161), 
        .B2(\completionDataOut[2][34] ), .ZN(n1952) );
  AOI22D1 U2418 ( .A1(n1175), .A2(\completionDataOut[1][33] ), .B1(n1187), 
        .B2(\completionDataOut[3][33] ), .ZN(n1949) );
  AOI22D1 U2419 ( .A1(n1150), .A2(\completionDataOut[0][33] ), .B1(n1161), 
        .B2(\completionDataOut[2][33] ), .ZN(n1948) );
  AOI22D1 U2420 ( .A1(n1175), .A2(\completionDataOut[1][32] ), .B1(n1187), 
        .B2(\completionDataOut[3][32] ), .ZN(n1945) );
  AOI22D1 U2421 ( .A1(n1150), .A2(\completionDataOut[0][32] ), .B1(n1161), 
        .B2(\completionDataOut[2][32] ), .ZN(n1944) );
  AOI22D1 U2422 ( .A1(n1226), .A2(\completionDataOut[5][31] ), .B1(n1237), 
        .B2(\completionDataOut[7][31] ), .ZN(n1943) );
  AOI22D1 U2423 ( .A1(n1201), .A2(\completionDataOut[4][31] ), .B1(n1212), 
        .B2(\completionDataOut[6][31] ), .ZN(n1942) );
  AOI22D1 U2424 ( .A1(n1175), .A2(\completionDataOut[1][31] ), .B1(n1187), 
        .B2(\completionDataOut[3][31] ), .ZN(n1941) );
  AOI22D1 U2425 ( .A1(n1150), .A2(\completionDataOut[0][31] ), .B1(n1161), 
        .B2(\completionDataOut[2][31] ), .ZN(n1940) );
  AOI22D1 U2426 ( .A1(n1226), .A2(\completionDataOut[5][30] ), .B1(n1237), 
        .B2(\completionDataOut[7][30] ), .ZN(n1939) );
  AOI22D1 U2427 ( .A1(n1201), .A2(\completionDataOut[4][30] ), .B1(n1212), 
        .B2(\completionDataOut[6][30] ), .ZN(n1938) );
  AOI22D1 U2428 ( .A1(n1175), .A2(\completionDataOut[1][30] ), .B1(n1187), 
        .B2(\completionDataOut[3][30] ), .ZN(n1937) );
  AOI22D1 U2429 ( .A1(n1150), .A2(\completionDataOut[0][30] ), .B1(n1161), 
        .B2(\completionDataOut[2][30] ), .ZN(n1936) );
  CKBD1 U2430 ( .I(n1245), .Z(n1237) );
  CKBD1 U2431 ( .I(n1231), .Z(n1226) );
  CKBD1 U2432 ( .I(n1220), .Z(n1212) );
  CKBD1 U2433 ( .I(n1206), .Z(n1201) );
  CKBD1 U2434 ( .I(n1180), .Z(n1175) );
  AOI22D1 U2435 ( .A1(n1150), .A2(\completionDataOut[0][29] ), .B1(n1161), 
        .B2(\completionDataOut[2][29] ), .ZN(n1935) );
  CKBD1 U2436 ( .I(n1169), .Z(n1161) );
  CKBD1 U2437 ( .I(n1155), .Z(n1150) );
  AOI22D1 U2438 ( .A1(n1231), .A2(\completionDataOut[5][24] ), .B1(n1238), 
        .B2(\completionDataOut[7][24] ), .ZN(n1918) );
  AOI22D1 U2439 ( .A1(n1206), .A2(\completionDataOut[4][24] ), .B1(n1213), 
        .B2(\completionDataOut[6][24] ), .ZN(n1917) );
  AOI22D1 U2440 ( .A1(n1180), .A2(\completionDataOut[1][24] ), .B1(n1188), 
        .B2(\completionDataOut[3][24] ), .ZN(n1916) );
  AOI22D1 U2441 ( .A1(n1155), .A2(\completionDataOut[0][24] ), .B1(n1162), 
        .B2(\completionDataOut[2][24] ), .ZN(n1915) );
  AOI22D1 U2442 ( .A1(n1155), .A2(\completionDataOut[0][23] ), .B1(n1162), 
        .B2(\completionDataOut[2][23] ), .ZN(n1914) );
  AOI22D1 U2443 ( .A1(n1176), .A2(\completionDataOut[1][22] ), .B1(n1189), 
        .B2(\completionDataOut[3][22] ), .ZN(n1911) );
  AOI22D1 U2444 ( .A1(n1151), .A2(\completionDataOut[0][22] ), .B1(n1163), 
        .B2(\completionDataOut[2][22] ), .ZN(n1910) );
  CKBD1 U2445 ( .I(n1241), .Z(n1239) );
  CKBD1 U2446 ( .I(n1230), .Z(n1227) );
  CKBD1 U2447 ( .I(n1233), .Z(n1230) );
  CKBD1 U2448 ( .I(n1216), .Z(n1214) );
  CKBD1 U2449 ( .I(n1205), .Z(n1202) );
  CKBD1 U2450 ( .I(n1208), .Z(n1205) );
  AOI22D1 U2451 ( .A1(n1176), .A2(\completionDataOut[1][21] ), .B1(n1189), 
        .B2(\completionDataOut[3][21] ), .ZN(n1907) );
  CKBD1 U2452 ( .I(n1191), .Z(n1189) );
  CKBD1 U2453 ( .I(n1179), .Z(n1176) );
  CKBD1 U2454 ( .I(n1182), .Z(n1179) );
  AOI22D1 U2455 ( .A1(n1151), .A2(\completionDataOut[0][21] ), .B1(n1163), 
        .B2(\completionDataOut[2][21] ), .ZN(n1906) );
  CKBD1 U2456 ( .I(n1165), .Z(n1163) );
  CKBD1 U2457 ( .I(n1169), .Z(n1165) );
  CKBD1 U2458 ( .I(n1154), .Z(n1151) );
  CKBD1 U2459 ( .I(n1157), .Z(n1154) );
  AOI22D1 U2460 ( .A1(n1180), .A2(\completionDataOut[1][27] ), .B1(n1188), 
        .B2(\completionDataOut[3][27] ), .ZN(n1928) );
  AOI22D1 U2461 ( .A1(n1155), .A2(\completionDataOut[0][27] ), .B1(n1162), 
        .B2(\completionDataOut[2][27] ), .ZN(n1927) );
  AOI22D1 U2462 ( .A1(n1180), .A2(\completionDataOut[1][26] ), .B1(n1188), 
        .B2(\completionDataOut[3][26] ), .ZN(n1924) );
  AOI22D1 U2463 ( .A1(n1155), .A2(\completionDataOut[0][26] ), .B1(n1162), 
        .B2(\completionDataOut[2][26] ), .ZN(n1923) );
  AOI22D1 U2464 ( .A1(n1231), .A2(\completionDataOut[5][25] ), .B1(n1238), 
        .B2(\completionDataOut[7][25] ), .ZN(n1922) );
  CKBD1 U2465 ( .I(n1246), .Z(n1238) );
  CKBD1 U2466 ( .I(n1233), .Z(n1231) );
  AOI22D1 U2467 ( .A1(n1206), .A2(\completionDataOut[4][25] ), .B1(n1213), 
        .B2(\completionDataOut[6][25] ), .ZN(n1921) );
  CKBD1 U2468 ( .I(n1221), .Z(n1213) );
  CKBD1 U2469 ( .I(n1208), .Z(n1206) );
  INVD1 U2470 ( .I(decodeReadAddr2_i[2]), .ZN(n2060) );
  AOI22D1 U2471 ( .A1(n1180), .A2(\completionDataOut[1][25] ), .B1(n1188), 
        .B2(\completionDataOut[3][25] ), .ZN(n1920) );
  NR2D1 U2472 ( .A1(decodeReadAddr2_i[2]), .A2(n1830), .ZN(n1831) );
  ND2D1 U2473 ( .A1(decodeReadAddr2_i[0]), .A2(decodeReadAddr2_i[1]), .ZN(
        n1830) );
  CKBD1 U2474 ( .I(n1182), .Z(n1180) );
  CKBD1 U2475 ( .I(n1183), .Z(n1182) );
  NR2D1 U2476 ( .A1(decodeReadAddr2_i[2]), .A2(n1828), .ZN(n1829) );
  INVD1 U2477 ( .I(decodeReadAddr2_i[1]), .ZN(n2059) );
  AOI22D1 U2478 ( .A1(n1155), .A2(\completionDataOut[0][25] ), .B1(n1162), 
        .B2(\completionDataOut[2][25] ), .ZN(n1919) );
  CKBD1 U2479 ( .I(n1170), .Z(n1162) );
  NR2D1 U2480 ( .A1(decodeReadAddr2_i[2]), .A2(n1826), .ZN(n1827) );
  ND2D1 U2481 ( .A1(decodeReadAddr2_i[1]), .A2(n2058), .ZN(n1826) );
  INVD1 U2482 ( .I(decodeReadAddr2_i[0]), .ZN(n2058) );
  CKBD1 U2483 ( .I(n1157), .Z(n1155) );
  AOI22D1 U2484 ( .A1(n1016), .A2(\completionDataOut[5][37] ), .B1(n1033), 
        .B2(\completionDataOut[7][37] ), .ZN(n1461) );
  CKBD1 U2485 ( .I(n1039), .Z(n1033) );
  NR2D1 U2486 ( .A1(n1592), .A2(n1308), .ZN(n1314) );
  AOI22D1 U2487 ( .A1(n984), .A2(\completionDataOut[4][37] ), .B1(n1001), .B2(
        \completionDataOut[6][37] ), .ZN(n1460) );
  CKBD1 U2488 ( .I(n1007), .Z(n1001) );
  CKBD1 U2489 ( .I(n996), .Z(n994) );
  CKBD1 U2490 ( .I(n1312), .Z(n996) );
  AOI22D1 U2491 ( .A1(n279), .A2(\completionDataOut[1][37] ), .B1(n969), .B2(
        \completionDataOut[3][37] ), .ZN(n1459) );
  CKBD1 U2492 ( .I(n975), .Z(n969) );
  AOI22D1 U2493 ( .A1(n288), .A2(\completionDataOut[0][37] ), .B1(n951), .B2(
        \completionDataOut[2][37] ), .ZN(n1458) );
  CKBD1 U2494 ( .I(n957), .Z(n951) );
  CKBD1 U2495 ( .I(n961), .Z(n957) );
  CKBD1 U2496 ( .I(n1305), .Z(n946) );
  CKBD1 U2497 ( .I(n938), .Z(n933) );
  CKBD1 U2498 ( .I(n885), .Z(n880) );
  CKBD1 U2499 ( .I(n819), .Z(n808) );
  CKBD1 U2500 ( .I(n915), .Z(n904) );
  CKBD1 U2501 ( .I(n914), .Z(n905) );
  CKBD1 U2502 ( .I(n940), .Z(n931) );
  CKBD1 U2503 ( .I(n942), .Z(n940) );
  CKBD1 U2504 ( .I(n941), .Z(n930) );
  CKBD1 U2505 ( .I(n942), .Z(n941) );
  CKBD1 U2506 ( .I(n899), .Z(n895) );
  CKBD1 U2507 ( .I(n899), .Z(n896) );
  CKBD1 U2508 ( .I(n901), .Z(n893) );
  CKBD1 U2509 ( .I(n901), .Z(n892) );
  CKBD1 U2510 ( .I(n913), .Z(n906) );
  CKBD1 U2511 ( .I(n888), .Z(n877) );
  CKBD1 U2512 ( .I(n889), .Z(n888) );
  CKBD1 U2513 ( .I(n887), .Z(n878) );
  CKBD1 U2514 ( .I(n889), .Z(n887) );
  CKBD1 U2515 ( .I(n819), .Z(n810) );
  CKBD1 U2516 ( .I(n819), .Z(n809) );
  CKBD1 U2517 ( .I(n821), .Z(n819) );
  CKBD1 U2518 ( .I(n828), .Z(n826) );
  CKBD1 U2519 ( .I(n834), .Z(n828) );
  CKBD1 U2520 ( .I(n829), .Z(n825) );
  CKBD1 U2521 ( .I(n834), .Z(n829) );
  CKBD1 U2522 ( .I(n858), .Z(n853) );
  CKBD1 U2523 ( .I(n900), .Z(n894) );
  CKBD1 U2524 ( .I(n912), .Z(n907) );
  CKBD1 U2525 ( .I(n898), .Z(n897) );
  CKBD1 U2526 ( .I(n910), .Z(n909) );
  CKBD1 U2527 ( .I(n927), .Z(n918) );
  CKBD1 U2528 ( .I(n927), .Z(n919) );
  CKBD1 U2529 ( .I(n939), .Z(n932) );
  CKBD1 U2530 ( .I(n942), .Z(n939) );
  CKBD1 U2531 ( .I(n925), .Z(n922) );
  CKBD1 U2532 ( .I(n937), .Z(n934) );
  CKBD1 U2533 ( .I(n925), .Z(n921) );
  CKBD1 U2534 ( .I(n871), .Z(n870) );
  CKBD1 U2535 ( .I(n883), .Z(n882) );
  CKBD1 U2536 ( .I(n873), .Z(n867) );
  INR2D1 U2537 ( .A1(n1303), .B1(n1302), .ZN(n2) );
  CKBD1 U2538 ( .I(n924), .Z(n923) );
  CKBD1 U2539 ( .I(n936), .Z(n935) );
  CKBD1 U2540 ( .I(n926), .Z(n920) );
  NR2D1 U2541 ( .A1(resets_i[7]), .A2(n1277), .ZN(n1280) );
  ND3D1 U2542 ( .A1(completionWriteAddr_i[0]), .A2(completionWriteAddr_i[1]), 
        .A3(n1278), .ZN(n1277) );
  CKBD1 U2543 ( .I(n872), .Z(n868) );
  CKBD1 U2544 ( .I(n884), .Z(n881) );
  CKBD1 U2545 ( .I(n874), .Z(n865) );
  CKBD1 U2546 ( .I(n886), .Z(n879) );
  CKBD1 U2547 ( .I(n872), .Z(n869) );
  CKBD1 U2548 ( .I(n874), .Z(n866) );
  CKBD1 U2549 ( .I(n889), .Z(n886) );
  NR2D1 U2550 ( .A1(resets_i[5]), .A2(n1270), .ZN(n1272) );
  ND2D1 U2551 ( .A1(n1278), .A2(n1303), .ZN(n1270) );
  CKBD1 U2552 ( .I(n844), .Z(n841) );
  CKBD1 U2553 ( .I(n857), .Z(n854) );
  CKBD1 U2554 ( .I(n846), .Z(n837) );
  CKBD1 U2555 ( .I(n844), .Z(n840) );
  CKBD1 U2556 ( .I(n843), .Z(n842) );
  CKBD1 U2557 ( .I(n856), .Z(n855) );
  CKBD1 U2558 ( .I(n845), .Z(n839) );
  CKBD1 U2559 ( .I(n846), .Z(n838) );
  CKBD1 U2560 ( .I(n859), .Z(n852) );
  CKBD1 U2561 ( .I(n862), .Z(n859) );
  CKBD1 U2562 ( .I(n861), .Z(n850) );
  CKBD1 U2563 ( .I(n862), .Z(n861) );
  CKBD1 U2564 ( .I(n860), .Z(n851) );
  CKBD1 U2565 ( .I(n862), .Z(n860) );
  NR2D1 U2566 ( .A1(resets_i[3]), .A2(n1266), .ZN(n1268) );
  IND3D1 U2567 ( .A1(n1302), .B1(completionWriteAddr_i[0]), .B2(
        completionWriteAddr_i[1]), .ZN(n1266) );
  CKBD1 U2568 ( .I(n817), .Z(n814) );
  CKBD1 U2569 ( .I(n831), .Z(n823) );
  CKBD1 U2570 ( .I(n833), .Z(n831) );
  CKBD1 U2571 ( .I(n818), .Z(n813) );
  CKBD1 U2572 ( .I(n830), .Z(n824) );
  CKBD1 U2573 ( .I(n833), .Z(n830) );
  CKBD1 U2574 ( .I(n832), .Z(n822) );
  CKBD1 U2575 ( .I(n833), .Z(n832) );
  CKBD1 U2576 ( .I(n816), .Z(n815) );
  NR2D1 U2577 ( .A1(resets_i[2]), .A2(n1263), .ZN(n1265) );
  INVD1 U2578 ( .I(completionWriteAddr_i[0]), .ZN(n1269) );
  NR2D1 U2579 ( .A1(n1299), .A2(n1291), .ZN(n1281) );
  ND2D1 U2580 ( .A1(decodeWriteAddr_i[1]), .A2(n1287), .ZN(n1291) );
  ND2D1 U2581 ( .A1(n1296), .A2(n1300), .ZN(n1288) );
  NR2D1 U2582 ( .A1(decodeWriteAddr_i[1]), .A2(n1287), .ZN(n1300) );
  INVD1 U2583 ( .I(decodeWriteAddr_i[0]), .ZN(n1287) );
  INVD1 U2584 ( .I(n1301), .ZN(n1296) );
  CKBD1 U2585 ( .I(n1027), .Z(n1025) );
  CKBD1 U2586 ( .I(n995), .Z(n993) );
  CKBD1 U2587 ( .I(n974), .Z(n980) );
  CKBD1 U2588 ( .I(n956), .Z(n962) );
  CKBD1 U2589 ( .I(n492), .Z(n1056) );
  CKBD1 U2590 ( .I(n1835), .Z(n1246) );
  CKBD1 U2591 ( .I(n1833), .Z(n1221) );
  CKBD1 U2592 ( .I(n493), .Z(n1157) );
  CKBD1 U2593 ( .I(n1314), .Z(n1028) );
  CKBD1 U2594 ( .I(n911), .Z(n908) );
  CKBD1 U2595 ( .I(n875), .Z(n872) );
  CKBD1 U2596 ( .I(n835), .Z(n834) );
  INR2D1 U2597 ( .A1(n1263), .B1(resets_i[2]), .ZN(n1264) );
  NR2D1 U2598 ( .A1(n1824), .A2(n1598), .ZN(n1603) );
  NR2D1 U2599 ( .A1(n1824), .A2(n1596), .ZN(n1602) );
  ND2D1 U2600 ( .A1(decodeReadAddr1_i[0]), .A2(n1823), .ZN(n1596) );
  NR2D1 U2601 ( .A1(n175), .A2(n1830), .ZN(n1835) );
  NR2D1 U2602 ( .A1(n175), .A2(n1826), .ZN(n1833) );
  ND2D1 U2603 ( .A1(decodeReadAddr2_i[0]), .A2(n2059), .ZN(n1828) );
  CKBD1 U2604 ( .I(n1315), .Z(n1043) );
  CKBD1 U2605 ( .I(n1313), .Z(n1011) );
  CKBD1 U2606 ( .I(n1311), .Z(n979) );
  CKBD1 U2607 ( .I(n1307), .Z(n961) );
  CKBD1 U2608 ( .I(n916), .Z(n915) );
  CKBD1 U2609 ( .I(n916), .Z(n914) );
  CKBD1 U2610 ( .I(n902), .Z(n899) );
  CKBD1 U2611 ( .I(n902), .Z(n901) );
  CKBD1 U2612 ( .I(n916), .Z(n913) );
  CKBD1 U2613 ( .I(n903), .Z(n900) );
  CKBD1 U2614 ( .I(n903), .Z(n898) );
  CKBD1 U2615 ( .I(n928), .Z(n927) );
  CKBD1 U2616 ( .I(n928), .Z(n925) );
  CKBD1 U2617 ( .I(n876), .Z(n871) );
  CKBD1 U2618 ( .I(n876), .Z(n873) );
  CKBD1 U2619 ( .I(n929), .Z(n924) );
  CKBD1 U2620 ( .I(n929), .Z(n926) );
  CKBD1 U2621 ( .I(n875), .Z(n874) );
  CKBD1 U2622 ( .I(n848), .Z(n843) );
  CKBD1 U2623 ( .I(n848), .Z(n845) );
  CKBD1 U2624 ( .I(n847), .Z(n846) );
  CKBD1 U2625 ( .I(n847), .Z(n844) );
  INR2D1 U2626 ( .A1(n1266), .B1(resets_i[3]), .ZN(n1267) );
  CKBD1 U2627 ( .I(n820), .Z(n817) );
  CKBD1 U2628 ( .I(n820), .Z(n818) );
  IND3D1 U2629 ( .A1(n1299), .B1(decodeWriteAddr_i[0]), .B2(
        decodeWriteAddr_i[1]), .ZN(n1284) );
  IND2D1 U2630 ( .A1(decodeWriteAddr_i[2]), .B1(decodeWriteEn_i), .ZN(n1299)
         );
  ND2D1 U2631 ( .A1(decodeWriteEn_i), .A2(decodeWriteAddr_i[2]), .ZN(n1301) );
  CKBD1 U2632 ( .I(n820), .Z(n816) );
  CKBD1 U2633 ( .I(n994), .Z(n987) );
  CKBD1 U2634 ( .I(n1026), .Z(n1019) );
  AO22D0 U2635 ( .A1(n835), .A2(\completionDataOut[2][6] ), .B1(n808), .B2(
        completionWriteData_i[6]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U2636 ( .A1(n835), .A2(\completionDataOut[2][7] ), .B1(n808), .B2(
        completionWriteData_i[7]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U2637 ( .A1(n835), .A2(\completionDataOut[2][8] ), .B1(n808), .B2(
        completionWriteData_i[8]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U2638 ( .A1(n835), .A2(\completionDataOut[2][9] ), .B1(n808), .B2(
        completionWriteData_i[9]), .Z(
        \eachCompletionReg[2].completionReg/eachEnDff[9].enDff/theFlop/N3 ) );
  AO22D0 U2639 ( .A1(n237), .A2(n863), .B1(n839), .B2(
        \completionDataOut[3][42] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[42].enDff/theFlop/N3 )
         );
  AO22D0 U2640 ( .A1(n248), .A2(n863), .B1(n840), .B2(
        \completionDataOut[3][53] ), .Z(
        \eachCompletionReg[3].completionReg/eachEnDff[53].enDff/theFlop/N3 )
         );
  AO22D0 U2641 ( .A1(completionWriteData_i[48]), .A2(n890), .B1(n867), .B2(
        \completionDataOut[5][48] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[48].enDff/theFlop/N3 )
         );
  AO22D0 U2642 ( .A1(completionWriteData_i[59]), .A2(n890), .B1(n869), .B2(
        \completionDataOut[5][59] ), .Z(
        \eachCompletionReg[5].completionReg/eachEnDff[59].enDff/theFlop/N3 )
         );
  AO22D0 U2643 ( .A1(n243), .A2(n494), .B1(n900), .B2(
        \completionDataOut[6][48] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[48].enDff/theFlop/N3 )
         );
  AO22D0 U2644 ( .A1(n254), .A2(n494), .B1(n896), .B2(
        \completionDataOut[6][59] ), .Z(
        \eachCompletionReg[6].completionReg/eachEnDff[59].enDff/theFlop/N3 )
         );
  AO22D0 U2645 ( .A1(n237), .A2(n943), .B1(n920), .B2(
        \completionDataOut[7][42] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[42].enDff/theFlop/N3 )
         );
  AO22D0 U2646 ( .A1(n248), .A2(n943), .B1(n921), .B2(
        \completionDataOut[7][53] ), .Z(
        \eachCompletionReg[7].completionReg/eachEnDff[53].enDff/theFlop/N3 )
         );
  AO22D0 U2647 ( .A1(n311), .A2(\managementDataOut[2][0] ), .B1(
        decodeWriteData_i[0]), .B2(n498), .Z(
        \eachManagementReg[2].managementReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U2648 ( .A1(n312), .A2(\managementDataOut[2][1] ), .B1(n498), .B2(
        decodeWriteData_i[1]), .Z(
        \eachManagementReg[2].managementReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U2649 ( .A1(n312), .A2(\managementDataOut[2][2] ), .B1(n498), .B2(
        decodeWriteData_i[2]), .Z(
        \eachManagementReg[2].managementReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U2650 ( .A1(n312), .A2(\managementDataOut[2][3] ), .B1(n498), .B2(
        decodeWriteData_i[3]), .Z(
        \eachManagementReg[2].managementReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U2651 ( .A1(n311), .A2(\managementDataOut[2][4] ), .B1(n499), .B2(
        decodeWriteData_i[4]), .Z(
        \eachManagementReg[2].managementReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U2652 ( .A1(n312), .A2(\managementDataOut[2][5] ), .B1(n499), .B2(
        decodeWriteData_i[5]), .Z(
        \eachManagementReg[2].managementReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U2653 ( .A1(n311), .A2(\managementDataOut[2][6] ), .B1(n499), .B2(
        decodeWriteData_i[6]), .Z(
        \eachManagementReg[2].managementReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U2654 ( .A1(n311), .A2(\managementDataOut[2][7] ), .B1(n499), .B2(
        decodeWriteData_i[7]), .Z(
        \eachManagementReg[2].managementReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U2655 ( .A1(n311), .A2(\managementDataOut[2][8] ), .B1(n499), .B2(
        decodeWriteData_i[8]), .Z(
        \eachManagementReg[2].managementReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U2656 ( .A1(n265), .A2(n506), .B1(n319), .B2(
        \managementDataOut[6][0] ), .Z(
        \eachManagementReg[6].managementReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U2657 ( .A1(n266), .A2(n506), .B1(n319), .B2(
        \managementDataOut[6][1] ), .Z(
        \eachManagementReg[6].managementReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U2658 ( .A1(n267), .A2(n506), .B1(n320), .B2(
        \managementDataOut[6][2] ), .Z(
        \eachManagementReg[6].managementReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U2659 ( .A1(n268), .A2(n506), .B1(n320), .B2(
        \managementDataOut[6][3] ), .Z(
        \eachManagementReg[6].managementReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U2660 ( .A1(n269), .A2(n506), .B1(n320), .B2(
        \managementDataOut[6][4] ), .Z(
        \eachManagementReg[6].managementReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U2661 ( .A1(n270), .A2(n507), .B1(n320), .B2(
        \managementDataOut[6][5] ), .Z(
        \eachManagementReg[6].managementReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U2662 ( .A1(n271), .A2(n507), .B1(n319), .B2(
        \managementDataOut[6][6] ), .Z(
        \eachManagementReg[6].managementReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U2663 ( .A1(n272), .A2(n507), .B1(n319), .B2(
        \managementDataOut[6][7] ), .Z(
        \eachManagementReg[6].managementReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U2664 ( .A1(n273), .A2(n507), .B1(n319), .B2(
        \managementDataOut[6][8] ), .Z(
        \eachManagementReg[6].managementReg/eachEnDff[8].enDff/theFlop/N3 ) );
endmodule


module ROB ( clk_i, reset_i, decodeReadAddr1_i, decodeReadAddr2_i, 
        decodeReadData1_o, decodeReadData2_o, updateTail_i, decodeWriteData_i, 
        nextTail_o, stall_o, completionWriteAddr_i, completionWriteEn_i, 
        completionWriteData_i, updateHead_i, head_o, commitReadData_o );
  input [3:0] decodeReadAddr1_i;
  input [3:0] decodeReadAddr2_i;
  output [64:0] decodeReadData1_o;
  output [64:0] decodeReadData2_o;
  input [8:0] decodeWriteData_i;
  output [3:0] nextTail_o;
  input [3:0] completionWriteAddr_i;
  input [69:0] completionWriteData_i;
  output [3:0] head_o;
  output [78:0] commitReadData_o;
  input clk_i, reset_i, updateTail_i, completionWriteEn_i, updateHead_i;
  output stall_o;
  wire   tailReset, decodeWriteEn, N6, N7, N8, N9, N10, N11, N12, N13,
         \headTailManager/headReset , \add_x_7/n1 , \add_x_6/n1 , n1, n3, n7,
         n11, n21, n25, n34, n35, n36, n37, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;
  wire   [2:0] tail;
  wire   [2:0] tailNext;
  wire   [2:0] head;
  wire   [2:0] decodeReadAddr1sub1;
  wire   [2:0] decodeReadAddr2sub1;
  wire   [2:0] completionWriteAddrsub1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9;
  assign head_o[3] = \add_x_7/n1 ;
  assign nextTail_o[3] = \add_x_6/n1 ;

  ROBregs theRegs ( .clk_i(clk_i), .resets_i({N13, n62, n64, n58, n61, n63, 
        n57, n59}), .decodeReadAddr1_i(decodeReadAddr1sub1), 
        .decodeReadAddr2_i(decodeReadAddr2sub1), .decodeWriteAddr_i({
        tailNext[2], n41, n48}), .decodeWriteEn_i(decodeWriteEn), 
        .decodeReadData1_o({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, decodeReadData1_o}), .decodeReadData2_o({
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, decodeReadData2_o}), .decodeWriteData_i(
        decodeWriteData_i), .completionWriteAddr_i(completionWriteAddrsub1), 
        .completionWriteEn_i(completionWriteEn_i), .completionWriteData_i(
        completionWriteData_i), .commitReadAddr_i({n51, head[1], n42}), 
        .commitReadData_o(commitReadData_o) );
  DFQD1 \headTailManager/headReset_reg  ( .D(n37), .CP(clk_i), .Q(
        \headTailManager/headReset ) );
  DFD1 \headTailManager/tail_reg[0]  ( .D(n34), .CP(clk_i), .Q(tail[0]), .QN(
        n65) );
  EDFKCND4 \headTailManager/head_reg[1]  ( .CN(n25), .D(head_o[1]), .E(
        updateHead_i), .CP(clk_i), .Q(head[1]), .QN(n40) );
  DFD2 \headTailManager/head_reg[0]  ( .D(n36), .CP(clk_i), .Q(head[0]), .QN(
        head_o[0]) );
  EDFKCND2 \headTailManager/tail_reg[1]  ( .CN(n21), .D(n1), .E(decodeWriteEn), 
        .CP(clk_i), .Q(tail[1]) );
  EDFKCND1 \headTailManager/head_reg[2]  ( .CN(n25), .D(head_o[2]), .E(
        updateHead_i), .CP(clk_i), .Q(n43), .QN(n50) );
  DFD2 \headTailManager/tailReset_reg  ( .D(n35), .CP(clk_i), .Q(tailReset), 
        .QN(n67) );
  EDFKCND2 \headTailManager/tail_reg[2]  ( .CN(n21), .D(n3), .E(decodeWriteEn), 
        .CP(clk_i), .Q(n66), .QN(n11) );
  CKND0 U52 ( .I(updateHead_i), .ZN(n60) );
  OA31D0 U53 ( .A1(n51), .A2(n71), .A3(n76), .B(n56), .Z(N8) );
  INVD2 U54 ( .I(N11), .ZN(n64) );
  XOR2D2 U55 ( .A1(decodeReadAddr1_i[2]), .A2(n68), .Z(decodeReadAddr1sub1[2])
         );
  ND2D1 U56 ( .A1(tail[0]), .A2(tail[1]), .ZN(n72) );
  NR2XD0 U57 ( .A1(n85), .A2(n84), .ZN(\add_x_6/n1 ) );
  INVD1 U58 ( .I(n46), .ZN(n41) );
  CKND2D2 U59 ( .A1(n42), .A2(n53), .ZN(n78) );
  CKND2 U60 ( .I(head_o[0]), .ZN(n42) );
  INVD2 U61 ( .I(n43), .ZN(n44) );
  INVD1 U62 ( .I(n40), .ZN(n53) );
  NR2XD0 U63 ( .A1(completionWriteAddr_i[1]), .A2(completionWriteAddr_i[0]), 
        .ZN(n70) );
  ND2D1 U64 ( .A1(n49), .A2(n47), .ZN(n84) );
  INVD1 U65 ( .I(N6), .ZN(n59) );
  INVD1 U66 ( .I(N10), .ZN(n58) );
  INVD1 U67 ( .I(N7), .ZN(n57) );
  AO21D1 U68 ( .A1(updateHead_i), .A2(\add_x_7/n1 ), .B(reset_i), .Z(N13) );
  OA31D1 U69 ( .A1(n44), .A2(n71), .A3(n76), .B(n55), .Z(N12) );
  OA31D1 U70 ( .A1(n44), .A2(n71), .A3(n77), .B(n56), .Z(N11) );
  CKBD1 U71 ( .I(n79), .Z(n54) );
  OA31D1 U72 ( .A1(n43), .A2(n71), .A3(n78), .B(n56), .Z(N9) );
  OA31D1 U73 ( .A1(n53), .A2(n43), .A3(n80), .B(n56), .Z(N6) );
  OA31D1 U74 ( .A1(n53), .A2(n44), .A3(n80), .B(n55), .Z(N10) );
  OA31D1 U75 ( .A1(n43), .A2(n71), .A3(n77), .B(n55), .Z(N7) );
  CKND2D0 U76 ( .A1(n77), .A2(n76), .ZN(head_o[1]) );
  OR2XD1 U77 ( .A1(n53), .A2(head_o[0]), .Z(n77) );
  INVD1 U78 ( .I(n60), .ZN(n45) );
  OAI21D1 U79 ( .A1(\headTailManager/headReset ), .A2(n81), .B(n56), .ZN(n79)
         );
  CKND1 U80 ( .I(n40), .ZN(n52) );
  INVD1 U81 ( .I(reset_i), .ZN(n55) );
  AO22D1 U82 ( .A1(tailReset), .A2(tail[0]), .B1(n65), .B2(n67), .Z(n7) );
  NR2XD0 U83 ( .A1(decodeReadAddr2_i[1]), .A2(decodeReadAddr2_i[0]), .ZN(n69)
         );
  NR2XD0 U84 ( .A1(decodeReadAddr1_i[1]), .A2(decodeReadAddr1_i[0]), .ZN(n68)
         );
  INVD1 U85 ( .I(tailNext[1]), .ZN(n46) );
  OA22D0 U86 ( .A1(n67), .A2(n1), .B1(tail[1]), .B2(tailReset), .Z(tailNext[1]) );
  INVD1 U87 ( .I(n46), .ZN(n47) );
  INVD1 U88 ( .I(n7), .ZN(n48) );
  INVD1 U89 ( .I(n7), .ZN(n49) );
  INVD1 U90 ( .I(n50), .ZN(n51) );
  AOI21D2 U91 ( .A1(n44), .A2(n78), .B(\add_x_7/n1 ), .ZN(head_o[2]) );
  ND2D1 U92 ( .A1(n52), .A2(head_o[0]), .ZN(n76) );
  INVD1 U93 ( .I(reset_i), .ZN(n56) );
  INVD1 U94 ( .I(n45), .ZN(n71) );
  AOI221D4 U95 ( .A1(updateTail_i), .A2(n83), .B1(n65), .B2(n83), .C(reset_i), 
        .ZN(n34) );
  AOI221D4 U96 ( .A1(n45), .A2(n80), .B1(head_o[0]), .B2(n80), .C(n54), .ZN(
        n36) );
  ND2D1 U97 ( .A1(n45), .A2(head_o[0]), .ZN(n80) );
  INVD1 U98 ( .I(decodeReadAddr1_i[0]), .ZN(decodeReadAddr1sub1[0]) );
  INVD1 U99 ( .I(decodeReadAddr2_i[0]), .ZN(decodeReadAddr2sub1[0]) );
  MUX2ND1 U100 ( .I0(n65), .I1(tail[0]), .S(tail[1]), .ZN(n1) );
  INVD1 U101 ( .I(N9), .ZN(n61) );
  OAI221D4 U102 ( .A1(n74), .A2(n53), .B1(n44), .B2(n3), .C(n73), .ZN(n75) );
  AOI22D2 U103 ( .A1(n52), .A2(n74), .B1(n3), .B2(n50), .ZN(n73) );
  OAI22D4 U104 ( .A1(n67), .A2(n3), .B1(n66), .B2(tailReset), .ZN(n85) );
  MUX2ND2 U105 ( .I0(n66), .I1(n11), .S(n72), .ZN(n3) );
  INVD1 U106 ( .I(N12), .ZN(n62) );
  INVD1 U107 ( .I(N8), .ZN(n63) );
  AOI21D2 U108 ( .A1(updateTail_i), .A2(n67), .B(reset_i), .ZN(n21) );
  AO21D2 U109 ( .A1(completionWriteAddr_i[0]), .A2(completionWriteAddr_i[1]), 
        .B(n70), .Z(completionWriteAddrsub1[1]) );
  AO21D1 U110 ( .A1(decodeReadAddr1_i[0]), .A2(decodeReadAddr1_i[1]), .B(n68), 
        .Z(decodeReadAddr1sub1[1]) );
  AO21D1 U111 ( .A1(decodeReadAddr2_i[0]), .A2(decodeReadAddr2_i[1]), .B(n69), 
        .Z(decodeReadAddr2sub1[1]) );
  NR2D2 U112 ( .A1(n44), .A2(n78), .ZN(\add_x_7/n1 ) );
  INVD1 U113 ( .I(completionWriteAddr_i[0]), .ZN(completionWriteAddrsub1[0])
         );
  OAI221D4 U114 ( .A1(tail[0]), .A2(decodeWriteEn), .B1(n65), .B2(n82), .C(
        tailReset), .ZN(n83) );
  NR2D3 U115 ( .A1(n82), .A2(n81), .ZN(decodeWriteEn) );
  AOI221D4 U116 ( .A1(tail[0]), .A2(head[0]), .B1(n65), .B2(head_o[0]), .C(n75), .ZN(n82) );
  OA21D1 U117 ( .A1(n49), .A2(n47), .B(n84), .Z(nextTail_o[1]) );
  INVD1 U118 ( .I(n49), .ZN(nextTail_o[0]) );
  CKXOR2D1 U119 ( .A1(decodeReadAddr2_i[2]), .A2(n69), .Z(
        decodeReadAddr2sub1[2]) );
  INVD1 U120 ( .I(n54), .ZN(n25) );
  CKXOR2D1 U121 ( .A1(completionWriteAddr_i[2]), .A2(n70), .Z(
        completionWriteAddrsub1[2]) );
  INVD1 U122 ( .I(n85), .ZN(tailNext[2]) );
  INVD1 U123 ( .I(updateTail_i), .ZN(n81) );
  INVD1 U124 ( .I(n1), .ZN(n74) );
  AOI21D1 U125 ( .A1(n85), .A2(n84), .B(\add_x_6/n1 ), .ZN(nextTail_o[2]) );
  INR2D1 U126 ( .A1(n82), .B1(n81), .ZN(stall_o) );
  AOI21D1 U127 ( .A1(n67), .A2(n81), .B(reset_i), .ZN(n35) );
  OA31D0 U128 ( .A1(updateTail_i), .A2(updateHead_i), .A3(
        \headTailManager/headReset ), .B(n56), .Z(n37) );
endmodule

