../../src/verilog/mux_4x1_X65.sv