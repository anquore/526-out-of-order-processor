library verilog;
use verilog.vl_types.all;
entity mux32x64_testbench is
end mux32x64_testbench;
