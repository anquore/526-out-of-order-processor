../../src/verilog/individualReg64.sv