library verilog;
use verilog.vl_types.all;
entity signExtend12_testbench is
end signExtend12_testbench;
