library verilog;
use verilog.vl_types.all;
entity andifier_testbench is
end andifier_testbench;
