../../src/verilog/wallOfDFFs.sv