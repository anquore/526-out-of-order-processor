../../src/verilog/dataMovement.sv