../../src/verilog/ALUStage.sv