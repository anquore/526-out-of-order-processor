library verilog;
use verilog.vl_types.all;
entity xnorifier_testbench is
end xnorifier_testbench;
