../../src/verilog/pipelinedProcessor.sv