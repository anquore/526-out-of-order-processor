../../src/verilog/decoder4x16.sv