../../src/verilog/completeDataPath.sv