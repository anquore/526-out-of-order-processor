../../src/verilog/fullReg32x64.sv