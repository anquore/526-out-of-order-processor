../../src/verilog/completeDataPathPipelined.sv