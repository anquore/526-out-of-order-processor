../../src/verilog/adderC65.sv