../../src/verilog/mapTable.sv