library verilog;
use verilog.vl_types.all;
entity mux8x1_testbench is
end mux8x1_testbench;
