../../src/verilog/mux2x5.sv