../../src/verilog/decoder2x4.sv