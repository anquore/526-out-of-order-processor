
module pipelined ( clk, reset );
  input clk, reset;


endmodule

