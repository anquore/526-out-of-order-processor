../../src/verilog/reservationStation.sv