../../src/verilog/reservationStationx2.sv