../../src/verilog/andifier.sv