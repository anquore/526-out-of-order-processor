library verilog;
use verilog.vl_types.all;
entity fullAdder_testbench is
end fullAdder_testbench;
