
module ROB ( clk_i, reset_i, decodeReadAddr1_i, decodeReadAddr2_i, 
        decodeReadData1_o, decodeReadData2_o, updateTail_i, decodeWriteData_i, 
        nextTail_o, stall_o, completionWriteAddr_i, completionWriteEn_i, 
        completionWriteData_i, updateHead_i, head_o, commitReadData_o );
  input [3:0] decodeReadAddr1_i;
  input [3:0] decodeReadAddr2_i;
  output [64:0] decodeReadData1_o;
  output [64:0] decodeReadData2_o;
  input [8:0] decodeWriteData_i;
  output [3:0] nextTail_o;
  input [3:0] completionWriteAddr_i;
  input [69:0] completionWriteData_i;
  output [3:0] head_o;
  output [78:0] commitReadData_o;
  input clk_i, reset_i, updateTail_i, completionWriteEn_i, updateHead_i;
  output stall_o;
  wire   n4118, tailReset, \headTailManager/headReset ,
         \theRegs/completionDataOut[0][0] , \theRegs/completionDataOut[0][1] ,
         \theRegs/completionDataOut[0][2] , \theRegs/completionDataOut[0][3] ,
         \theRegs/completionDataOut[0][4] , \theRegs/completionDataOut[0][5] ,
         \theRegs/completionDataOut[0][6] , \theRegs/completionDataOut[0][7] ,
         \theRegs/completionDataOut[0][8] , \theRegs/completionDataOut[0][9] ,
         \theRegs/completionDataOut[0][10] ,
         \theRegs/completionDataOut[0][11] ,
         \theRegs/completionDataOut[0][12] ,
         \theRegs/completionDataOut[0][13] ,
         \theRegs/completionDataOut[0][14] ,
         \theRegs/completionDataOut[0][15] ,
         \theRegs/completionDataOut[0][16] ,
         \theRegs/completionDataOut[0][17] ,
         \theRegs/completionDataOut[0][18] ,
         \theRegs/completionDataOut[0][19] ,
         \theRegs/completionDataOut[0][20] ,
         \theRegs/completionDataOut[0][21] ,
         \theRegs/completionDataOut[0][22] ,
         \theRegs/completionDataOut[0][23] ,
         \theRegs/completionDataOut[0][24] ,
         \theRegs/completionDataOut[0][25] ,
         \theRegs/completionDataOut[0][26] ,
         \theRegs/completionDataOut[0][27] ,
         \theRegs/completionDataOut[0][28] ,
         \theRegs/completionDataOut[0][29] ,
         \theRegs/completionDataOut[0][30] ,
         \theRegs/completionDataOut[0][31] ,
         \theRegs/completionDataOut[0][32] ,
         \theRegs/completionDataOut[0][33] ,
         \theRegs/completionDataOut[0][34] ,
         \theRegs/completionDataOut[0][35] ,
         \theRegs/completionDataOut[0][36] ,
         \theRegs/completionDataOut[0][37] ,
         \theRegs/completionDataOut[0][38] ,
         \theRegs/completionDataOut[0][39] ,
         \theRegs/completionDataOut[0][40] ,
         \theRegs/completionDataOut[0][41] ,
         \theRegs/completionDataOut[0][42] ,
         \theRegs/completionDataOut[0][43] ,
         \theRegs/completionDataOut[0][44] ,
         \theRegs/completionDataOut[0][45] ,
         \theRegs/completionDataOut[0][46] ,
         \theRegs/completionDataOut[0][47] ,
         \theRegs/completionDataOut[0][48] ,
         \theRegs/completionDataOut[0][49] ,
         \theRegs/completionDataOut[0][50] ,
         \theRegs/completionDataOut[0][51] ,
         \theRegs/completionDataOut[0][52] ,
         \theRegs/completionDataOut[0][53] ,
         \theRegs/completionDataOut[0][54] ,
         \theRegs/completionDataOut[0][55] ,
         \theRegs/completionDataOut[0][56] ,
         \theRegs/completionDataOut[0][57] ,
         \theRegs/completionDataOut[0][58] ,
         \theRegs/completionDataOut[0][59] ,
         \theRegs/completionDataOut[0][60] ,
         \theRegs/completionDataOut[0][61] ,
         \theRegs/completionDataOut[0][62] ,
         \theRegs/completionDataOut[0][63] ,
         \theRegs/completionDataOut[0][64] ,
         \theRegs/completionDataOut[0][65] ,
         \theRegs/completionDataOut[0][66] ,
         \theRegs/completionDataOut[0][67] ,
         \theRegs/completionDataOut[0][68] ,
         \theRegs/completionDataOut[0][69] , \theRegs/completionDataOut[1][0] ,
         \theRegs/completionDataOut[1][1] , \theRegs/completionDataOut[1][2] ,
         \theRegs/completionDataOut[1][3] , \theRegs/completionDataOut[1][4] ,
         \theRegs/completionDataOut[1][5] , \theRegs/completionDataOut[1][6] ,
         \theRegs/completionDataOut[1][7] , \theRegs/completionDataOut[1][8] ,
         \theRegs/completionDataOut[1][9] , \theRegs/completionDataOut[1][10] ,
         \theRegs/completionDataOut[1][11] ,
         \theRegs/completionDataOut[1][12] ,
         \theRegs/completionDataOut[1][13] ,
         \theRegs/completionDataOut[1][14] ,
         \theRegs/completionDataOut[1][15] ,
         \theRegs/completionDataOut[1][16] ,
         \theRegs/completionDataOut[1][17] ,
         \theRegs/completionDataOut[1][18] ,
         \theRegs/completionDataOut[1][19] ,
         \theRegs/completionDataOut[1][20] ,
         \theRegs/completionDataOut[1][21] ,
         \theRegs/completionDataOut[1][22] ,
         \theRegs/completionDataOut[1][23] ,
         \theRegs/completionDataOut[1][24] ,
         \theRegs/completionDataOut[1][25] ,
         \theRegs/completionDataOut[1][26] ,
         \theRegs/completionDataOut[1][27] ,
         \theRegs/completionDataOut[1][28] ,
         \theRegs/completionDataOut[1][29] ,
         \theRegs/completionDataOut[1][30] ,
         \theRegs/completionDataOut[1][31] ,
         \theRegs/completionDataOut[1][32] ,
         \theRegs/completionDataOut[1][33] ,
         \theRegs/completionDataOut[1][34] ,
         \theRegs/completionDataOut[1][35] ,
         \theRegs/completionDataOut[1][36] ,
         \theRegs/completionDataOut[1][37] ,
         \theRegs/completionDataOut[1][38] ,
         \theRegs/completionDataOut[1][39] ,
         \theRegs/completionDataOut[1][40] ,
         \theRegs/completionDataOut[1][41] ,
         \theRegs/completionDataOut[1][42] ,
         \theRegs/completionDataOut[1][43] ,
         \theRegs/completionDataOut[1][44] ,
         \theRegs/completionDataOut[1][45] ,
         \theRegs/completionDataOut[1][46] ,
         \theRegs/completionDataOut[1][47] ,
         \theRegs/completionDataOut[1][48] ,
         \theRegs/completionDataOut[1][49] ,
         \theRegs/completionDataOut[1][50] ,
         \theRegs/completionDataOut[1][51] ,
         \theRegs/completionDataOut[1][52] ,
         \theRegs/completionDataOut[1][53] ,
         \theRegs/completionDataOut[1][54] ,
         \theRegs/completionDataOut[1][55] ,
         \theRegs/completionDataOut[1][56] ,
         \theRegs/completionDataOut[1][57] ,
         \theRegs/completionDataOut[1][58] ,
         \theRegs/completionDataOut[1][59] ,
         \theRegs/completionDataOut[1][60] ,
         \theRegs/completionDataOut[1][61] ,
         \theRegs/completionDataOut[1][62] ,
         \theRegs/completionDataOut[1][63] ,
         \theRegs/completionDataOut[1][64] ,
         \theRegs/completionDataOut[1][65] ,
         \theRegs/completionDataOut[1][66] ,
         \theRegs/completionDataOut[1][67] ,
         \theRegs/completionDataOut[1][68] ,
         \theRegs/completionDataOut[1][69] , \theRegs/completionDataOut[2][0] ,
         \theRegs/completionDataOut[2][1] , \theRegs/completionDataOut[2][2] ,
         \theRegs/completionDataOut[2][3] , \theRegs/completionDataOut[2][4] ,
         \theRegs/completionDataOut[2][5] , \theRegs/completionDataOut[2][6] ,
         \theRegs/completionDataOut[2][7] , \theRegs/completionDataOut[2][8] ,
         \theRegs/completionDataOut[2][9] , \theRegs/completionDataOut[2][10] ,
         \theRegs/completionDataOut[2][11] ,
         \theRegs/completionDataOut[2][12] ,
         \theRegs/completionDataOut[2][13] ,
         \theRegs/completionDataOut[2][14] ,
         \theRegs/completionDataOut[2][15] ,
         \theRegs/completionDataOut[2][16] ,
         \theRegs/completionDataOut[2][17] ,
         \theRegs/completionDataOut[2][18] ,
         \theRegs/completionDataOut[2][19] ,
         \theRegs/completionDataOut[2][20] ,
         \theRegs/completionDataOut[2][21] ,
         \theRegs/completionDataOut[2][22] ,
         \theRegs/completionDataOut[2][23] ,
         \theRegs/completionDataOut[2][24] ,
         \theRegs/completionDataOut[2][25] ,
         \theRegs/completionDataOut[2][26] ,
         \theRegs/completionDataOut[2][27] ,
         \theRegs/completionDataOut[2][28] ,
         \theRegs/completionDataOut[2][29] ,
         \theRegs/completionDataOut[2][30] ,
         \theRegs/completionDataOut[2][31] ,
         \theRegs/completionDataOut[2][32] ,
         \theRegs/completionDataOut[2][33] ,
         \theRegs/completionDataOut[2][34] ,
         \theRegs/completionDataOut[2][35] ,
         \theRegs/completionDataOut[2][36] ,
         \theRegs/completionDataOut[2][37] ,
         \theRegs/completionDataOut[2][38] ,
         \theRegs/completionDataOut[2][39] ,
         \theRegs/completionDataOut[2][40] ,
         \theRegs/completionDataOut[2][41] ,
         \theRegs/completionDataOut[2][42] ,
         \theRegs/completionDataOut[2][43] ,
         \theRegs/completionDataOut[2][44] ,
         \theRegs/completionDataOut[2][45] ,
         \theRegs/completionDataOut[2][46] ,
         \theRegs/completionDataOut[2][47] ,
         \theRegs/completionDataOut[2][48] ,
         \theRegs/completionDataOut[2][49] ,
         \theRegs/completionDataOut[2][50] ,
         \theRegs/completionDataOut[2][51] ,
         \theRegs/completionDataOut[2][52] ,
         \theRegs/completionDataOut[2][53] ,
         \theRegs/completionDataOut[2][54] ,
         \theRegs/completionDataOut[2][55] ,
         \theRegs/completionDataOut[2][56] ,
         \theRegs/completionDataOut[2][57] ,
         \theRegs/completionDataOut[2][58] ,
         \theRegs/completionDataOut[2][59] ,
         \theRegs/completionDataOut[2][60] ,
         \theRegs/completionDataOut[2][61] ,
         \theRegs/completionDataOut[2][62] ,
         \theRegs/completionDataOut[2][63] ,
         \theRegs/completionDataOut[2][64] ,
         \theRegs/completionDataOut[2][65] ,
         \theRegs/completionDataOut[2][66] ,
         \theRegs/completionDataOut[2][67] ,
         \theRegs/completionDataOut[2][68] ,
         \theRegs/completionDataOut[2][69] , \theRegs/completionDataOut[3][0] ,
         \theRegs/completionDataOut[3][1] , \theRegs/completionDataOut[3][2] ,
         \theRegs/completionDataOut[3][3] , \theRegs/completionDataOut[3][4] ,
         \theRegs/completionDataOut[3][5] , \theRegs/completionDataOut[3][6] ,
         \theRegs/completionDataOut[3][7] , \theRegs/completionDataOut[3][8] ,
         \theRegs/completionDataOut[3][9] , \theRegs/completionDataOut[3][10] ,
         \theRegs/completionDataOut[3][11] ,
         \theRegs/completionDataOut[3][12] ,
         \theRegs/completionDataOut[3][13] ,
         \theRegs/completionDataOut[3][14] ,
         \theRegs/completionDataOut[3][15] ,
         \theRegs/completionDataOut[3][16] ,
         \theRegs/completionDataOut[3][17] ,
         \theRegs/completionDataOut[3][18] ,
         \theRegs/completionDataOut[3][19] ,
         \theRegs/completionDataOut[3][20] ,
         \theRegs/completionDataOut[3][21] ,
         \theRegs/completionDataOut[3][22] ,
         \theRegs/completionDataOut[3][23] ,
         \theRegs/completionDataOut[3][24] ,
         \theRegs/completionDataOut[3][25] ,
         \theRegs/completionDataOut[3][26] ,
         \theRegs/completionDataOut[3][27] ,
         \theRegs/completionDataOut[3][28] ,
         \theRegs/completionDataOut[3][29] ,
         \theRegs/completionDataOut[3][30] ,
         \theRegs/completionDataOut[3][31] ,
         \theRegs/completionDataOut[3][32] ,
         \theRegs/completionDataOut[3][33] ,
         \theRegs/completionDataOut[3][34] ,
         \theRegs/completionDataOut[3][35] ,
         \theRegs/completionDataOut[3][36] ,
         \theRegs/completionDataOut[3][37] ,
         \theRegs/completionDataOut[3][38] ,
         \theRegs/completionDataOut[3][39] ,
         \theRegs/completionDataOut[3][40] ,
         \theRegs/completionDataOut[3][41] ,
         \theRegs/completionDataOut[3][42] ,
         \theRegs/completionDataOut[3][43] ,
         \theRegs/completionDataOut[3][44] ,
         \theRegs/completionDataOut[3][45] ,
         \theRegs/completionDataOut[3][46] ,
         \theRegs/completionDataOut[3][47] ,
         \theRegs/completionDataOut[3][48] ,
         \theRegs/completionDataOut[3][49] ,
         \theRegs/completionDataOut[3][50] ,
         \theRegs/completionDataOut[3][51] ,
         \theRegs/completionDataOut[3][52] ,
         \theRegs/completionDataOut[3][53] ,
         \theRegs/completionDataOut[3][54] ,
         \theRegs/completionDataOut[3][55] ,
         \theRegs/completionDataOut[3][56] ,
         \theRegs/completionDataOut[3][57] ,
         \theRegs/completionDataOut[3][58] ,
         \theRegs/completionDataOut[3][59] ,
         \theRegs/completionDataOut[3][60] ,
         \theRegs/completionDataOut[3][61] ,
         \theRegs/completionDataOut[3][62] ,
         \theRegs/completionDataOut[3][63] ,
         \theRegs/completionDataOut[3][64] ,
         \theRegs/completionDataOut[3][65] ,
         \theRegs/completionDataOut[3][66] ,
         \theRegs/completionDataOut[3][67] ,
         \theRegs/completionDataOut[3][68] ,
         \theRegs/completionDataOut[3][69] , \theRegs/completionDataOut[4][0] ,
         \theRegs/completionDataOut[4][1] , \theRegs/completionDataOut[4][2] ,
         \theRegs/completionDataOut[4][3] , \theRegs/completionDataOut[4][4] ,
         \theRegs/completionDataOut[4][5] , \theRegs/completionDataOut[4][6] ,
         \theRegs/completionDataOut[4][7] , \theRegs/completionDataOut[4][8] ,
         \theRegs/completionDataOut[4][9] , \theRegs/completionDataOut[4][10] ,
         \theRegs/completionDataOut[4][11] ,
         \theRegs/completionDataOut[4][12] ,
         \theRegs/completionDataOut[4][13] ,
         \theRegs/completionDataOut[4][14] ,
         \theRegs/completionDataOut[4][15] ,
         \theRegs/completionDataOut[4][16] ,
         \theRegs/completionDataOut[4][17] ,
         \theRegs/completionDataOut[4][18] ,
         \theRegs/completionDataOut[4][19] ,
         \theRegs/completionDataOut[4][20] ,
         \theRegs/completionDataOut[4][21] ,
         \theRegs/completionDataOut[4][22] ,
         \theRegs/completionDataOut[4][23] ,
         \theRegs/completionDataOut[4][24] ,
         \theRegs/completionDataOut[4][25] ,
         \theRegs/completionDataOut[4][26] ,
         \theRegs/completionDataOut[4][27] ,
         \theRegs/completionDataOut[4][28] ,
         \theRegs/completionDataOut[4][29] ,
         \theRegs/completionDataOut[4][30] ,
         \theRegs/completionDataOut[4][31] ,
         \theRegs/completionDataOut[4][32] ,
         \theRegs/completionDataOut[4][33] ,
         \theRegs/completionDataOut[4][34] ,
         \theRegs/completionDataOut[4][35] ,
         \theRegs/completionDataOut[4][36] ,
         \theRegs/completionDataOut[4][37] ,
         \theRegs/completionDataOut[4][38] ,
         \theRegs/completionDataOut[4][39] ,
         \theRegs/completionDataOut[4][40] ,
         \theRegs/completionDataOut[4][41] ,
         \theRegs/completionDataOut[4][42] ,
         \theRegs/completionDataOut[4][43] ,
         \theRegs/completionDataOut[4][44] ,
         \theRegs/completionDataOut[4][45] ,
         \theRegs/completionDataOut[4][46] ,
         \theRegs/completionDataOut[4][47] ,
         \theRegs/completionDataOut[4][48] ,
         \theRegs/completionDataOut[4][49] ,
         \theRegs/completionDataOut[4][50] ,
         \theRegs/completionDataOut[4][51] ,
         \theRegs/completionDataOut[4][52] ,
         \theRegs/completionDataOut[4][53] ,
         \theRegs/completionDataOut[4][54] ,
         \theRegs/completionDataOut[4][55] ,
         \theRegs/completionDataOut[4][56] ,
         \theRegs/completionDataOut[4][57] ,
         \theRegs/completionDataOut[4][58] ,
         \theRegs/completionDataOut[4][59] ,
         \theRegs/completionDataOut[4][60] ,
         \theRegs/completionDataOut[4][61] ,
         \theRegs/completionDataOut[4][62] ,
         \theRegs/completionDataOut[4][63] ,
         \theRegs/completionDataOut[4][64] ,
         \theRegs/completionDataOut[4][65] ,
         \theRegs/completionDataOut[4][66] ,
         \theRegs/completionDataOut[4][67] ,
         \theRegs/completionDataOut[4][68] ,
         \theRegs/completionDataOut[4][69] , \theRegs/completionDataOut[5][0] ,
         \theRegs/completionDataOut[5][1] , \theRegs/completionDataOut[5][2] ,
         \theRegs/completionDataOut[5][3] , \theRegs/completionDataOut[5][4] ,
         \theRegs/completionDataOut[5][5] , \theRegs/completionDataOut[5][6] ,
         \theRegs/completionDataOut[5][7] , \theRegs/completionDataOut[5][8] ,
         \theRegs/completionDataOut[5][9] , \theRegs/completionDataOut[5][10] ,
         \theRegs/completionDataOut[5][11] ,
         \theRegs/completionDataOut[5][12] ,
         \theRegs/completionDataOut[5][13] ,
         \theRegs/completionDataOut[5][14] ,
         \theRegs/completionDataOut[5][15] ,
         \theRegs/completionDataOut[5][16] ,
         \theRegs/completionDataOut[5][17] ,
         \theRegs/completionDataOut[5][18] ,
         \theRegs/completionDataOut[5][19] ,
         \theRegs/completionDataOut[5][20] ,
         \theRegs/completionDataOut[5][21] ,
         \theRegs/completionDataOut[5][22] ,
         \theRegs/completionDataOut[5][23] ,
         \theRegs/completionDataOut[5][24] ,
         \theRegs/completionDataOut[5][25] ,
         \theRegs/completionDataOut[5][26] ,
         \theRegs/completionDataOut[5][27] ,
         \theRegs/completionDataOut[5][28] ,
         \theRegs/completionDataOut[5][29] ,
         \theRegs/completionDataOut[5][30] ,
         \theRegs/completionDataOut[5][31] ,
         \theRegs/completionDataOut[5][32] ,
         \theRegs/completionDataOut[5][33] ,
         \theRegs/completionDataOut[5][34] ,
         \theRegs/completionDataOut[5][35] ,
         \theRegs/completionDataOut[5][36] ,
         \theRegs/completionDataOut[5][37] ,
         \theRegs/completionDataOut[5][38] ,
         \theRegs/completionDataOut[5][39] ,
         \theRegs/completionDataOut[5][40] ,
         \theRegs/completionDataOut[5][41] ,
         \theRegs/completionDataOut[5][42] ,
         \theRegs/completionDataOut[5][43] ,
         \theRegs/completionDataOut[5][44] ,
         \theRegs/completionDataOut[5][45] ,
         \theRegs/completionDataOut[5][46] ,
         \theRegs/completionDataOut[5][47] ,
         \theRegs/completionDataOut[5][48] ,
         \theRegs/completionDataOut[5][49] ,
         \theRegs/completionDataOut[5][50] ,
         \theRegs/completionDataOut[5][51] ,
         \theRegs/completionDataOut[5][52] ,
         \theRegs/completionDataOut[5][53] ,
         \theRegs/completionDataOut[5][54] ,
         \theRegs/completionDataOut[5][55] ,
         \theRegs/completionDataOut[5][56] ,
         \theRegs/completionDataOut[5][57] ,
         \theRegs/completionDataOut[5][58] ,
         \theRegs/completionDataOut[5][59] ,
         \theRegs/completionDataOut[5][60] ,
         \theRegs/completionDataOut[5][61] ,
         \theRegs/completionDataOut[5][62] ,
         \theRegs/completionDataOut[5][63] ,
         \theRegs/completionDataOut[5][64] ,
         \theRegs/completionDataOut[5][65] ,
         \theRegs/completionDataOut[5][66] ,
         \theRegs/completionDataOut[5][67] ,
         \theRegs/completionDataOut[5][68] ,
         \theRegs/completionDataOut[5][69] , \theRegs/completionDataOut[6][0] ,
         \theRegs/completionDataOut[6][1] , \theRegs/completionDataOut[6][2] ,
         \theRegs/completionDataOut[6][3] , \theRegs/completionDataOut[6][4] ,
         \theRegs/completionDataOut[6][5] , \theRegs/completionDataOut[6][6] ,
         \theRegs/completionDataOut[6][7] , \theRegs/completionDataOut[6][8] ,
         \theRegs/completionDataOut[6][9] , \theRegs/completionDataOut[6][10] ,
         \theRegs/completionDataOut[6][11] ,
         \theRegs/completionDataOut[6][12] ,
         \theRegs/completionDataOut[6][13] ,
         \theRegs/completionDataOut[6][14] ,
         \theRegs/completionDataOut[6][15] ,
         \theRegs/completionDataOut[6][16] ,
         \theRegs/completionDataOut[6][17] ,
         \theRegs/completionDataOut[6][18] ,
         \theRegs/completionDataOut[6][19] ,
         \theRegs/completionDataOut[6][20] ,
         \theRegs/completionDataOut[6][21] ,
         \theRegs/completionDataOut[6][22] ,
         \theRegs/completionDataOut[6][23] ,
         \theRegs/completionDataOut[6][24] ,
         \theRegs/completionDataOut[6][25] ,
         \theRegs/completionDataOut[6][26] ,
         \theRegs/completionDataOut[6][27] ,
         \theRegs/completionDataOut[6][28] ,
         \theRegs/completionDataOut[6][29] ,
         \theRegs/completionDataOut[6][30] ,
         \theRegs/completionDataOut[6][31] ,
         \theRegs/completionDataOut[6][32] ,
         \theRegs/completionDataOut[6][33] ,
         \theRegs/completionDataOut[6][34] ,
         \theRegs/completionDataOut[6][35] ,
         \theRegs/completionDataOut[6][36] ,
         \theRegs/completionDataOut[6][37] ,
         \theRegs/completionDataOut[6][38] ,
         \theRegs/completionDataOut[6][39] ,
         \theRegs/completionDataOut[6][40] ,
         \theRegs/completionDataOut[6][41] ,
         \theRegs/completionDataOut[6][42] ,
         \theRegs/completionDataOut[6][43] ,
         \theRegs/completionDataOut[6][44] ,
         \theRegs/completionDataOut[6][45] ,
         \theRegs/completionDataOut[6][46] ,
         \theRegs/completionDataOut[6][47] ,
         \theRegs/completionDataOut[6][48] ,
         \theRegs/completionDataOut[6][49] ,
         \theRegs/completionDataOut[6][50] ,
         \theRegs/completionDataOut[6][51] ,
         \theRegs/completionDataOut[6][52] ,
         \theRegs/completionDataOut[6][53] ,
         \theRegs/completionDataOut[6][54] ,
         \theRegs/completionDataOut[6][55] ,
         \theRegs/completionDataOut[6][56] ,
         \theRegs/completionDataOut[6][57] ,
         \theRegs/completionDataOut[6][58] ,
         \theRegs/completionDataOut[6][59] ,
         \theRegs/completionDataOut[6][60] ,
         \theRegs/completionDataOut[6][61] ,
         \theRegs/completionDataOut[6][62] ,
         \theRegs/completionDataOut[6][63] ,
         \theRegs/completionDataOut[6][64] ,
         \theRegs/completionDataOut[6][65] ,
         \theRegs/completionDataOut[6][66] ,
         \theRegs/completionDataOut[6][67] ,
         \theRegs/completionDataOut[6][68] ,
         \theRegs/completionDataOut[6][69] , \theRegs/completionDataOut[7][0] ,
         \theRegs/completionDataOut[7][1] , \theRegs/completionDataOut[7][2] ,
         \theRegs/completionDataOut[7][3] , \theRegs/completionDataOut[7][4] ,
         \theRegs/completionDataOut[7][5] , \theRegs/completionDataOut[7][6] ,
         \theRegs/completionDataOut[7][7] , \theRegs/completionDataOut[7][8] ,
         \theRegs/completionDataOut[7][9] , \theRegs/completionDataOut[7][10] ,
         \theRegs/completionDataOut[7][11] ,
         \theRegs/completionDataOut[7][12] ,
         \theRegs/completionDataOut[7][13] ,
         \theRegs/completionDataOut[7][14] ,
         \theRegs/completionDataOut[7][15] ,
         \theRegs/completionDataOut[7][16] ,
         \theRegs/completionDataOut[7][17] ,
         \theRegs/completionDataOut[7][18] ,
         \theRegs/completionDataOut[7][19] ,
         \theRegs/completionDataOut[7][20] ,
         \theRegs/completionDataOut[7][21] ,
         \theRegs/completionDataOut[7][22] ,
         \theRegs/completionDataOut[7][23] ,
         \theRegs/completionDataOut[7][24] ,
         \theRegs/completionDataOut[7][25] ,
         \theRegs/completionDataOut[7][26] ,
         \theRegs/completionDataOut[7][27] ,
         \theRegs/completionDataOut[7][28] ,
         \theRegs/completionDataOut[7][29] ,
         \theRegs/completionDataOut[7][30] ,
         \theRegs/completionDataOut[7][31] ,
         \theRegs/completionDataOut[7][32] ,
         \theRegs/completionDataOut[7][33] ,
         \theRegs/completionDataOut[7][34] ,
         \theRegs/completionDataOut[7][35] ,
         \theRegs/completionDataOut[7][36] ,
         \theRegs/completionDataOut[7][37] ,
         \theRegs/completionDataOut[7][38] ,
         \theRegs/completionDataOut[7][39] ,
         \theRegs/completionDataOut[7][40] ,
         \theRegs/completionDataOut[7][41] ,
         \theRegs/completionDataOut[7][42] ,
         \theRegs/completionDataOut[7][43] ,
         \theRegs/completionDataOut[7][44] ,
         \theRegs/completionDataOut[7][45] ,
         \theRegs/completionDataOut[7][46] ,
         \theRegs/completionDataOut[7][47] ,
         \theRegs/completionDataOut[7][48] ,
         \theRegs/completionDataOut[7][49] ,
         \theRegs/completionDataOut[7][50] ,
         \theRegs/completionDataOut[7][51] ,
         \theRegs/completionDataOut[7][52] ,
         \theRegs/completionDataOut[7][53] ,
         \theRegs/completionDataOut[7][54] ,
         \theRegs/completionDataOut[7][55] ,
         \theRegs/completionDataOut[7][56] ,
         \theRegs/completionDataOut[7][57] ,
         \theRegs/completionDataOut[7][58] ,
         \theRegs/completionDataOut[7][59] ,
         \theRegs/completionDataOut[7][60] ,
         \theRegs/completionDataOut[7][61] ,
         \theRegs/completionDataOut[7][62] ,
         \theRegs/completionDataOut[7][63] ,
         \theRegs/completionDataOut[7][64] ,
         \theRegs/completionDataOut[7][65] ,
         \theRegs/completionDataOut[7][66] ,
         \theRegs/completionDataOut[7][67] ,
         \theRegs/completionDataOut[7][68] ,
         \theRegs/completionDataOut[7][69] , \theRegs/managementDataOut[7][8] ,
         \theRegs/managementDataOut[7][7] , \theRegs/managementDataOut[7][6] ,
         \theRegs/managementDataOut[7][5] , \theRegs/managementDataOut[7][4] ,
         \theRegs/managementDataOut[7][3] , \theRegs/managementDataOut[7][2] ,
         \theRegs/managementDataOut[7][1] , \theRegs/managementDataOut[7][0] ,
         \theRegs/managementDataOut[6][8] , \theRegs/managementDataOut[6][7] ,
         \theRegs/managementDataOut[6][6] , \theRegs/managementDataOut[6][5] ,
         \theRegs/managementDataOut[6][4] , \theRegs/managementDataOut[6][3] ,
         \theRegs/managementDataOut[6][2] , \theRegs/managementDataOut[6][1] ,
         \theRegs/managementDataOut[6][0] , \theRegs/managementDataOut[5][8] ,
         \theRegs/managementDataOut[5][7] , \theRegs/managementDataOut[5][6] ,
         \theRegs/managementDataOut[5][5] , \theRegs/managementDataOut[5][4] ,
         \theRegs/managementDataOut[5][3] , \theRegs/managementDataOut[5][2] ,
         \theRegs/managementDataOut[5][1] , \theRegs/managementDataOut[5][0] ,
         \theRegs/managementDataOut[4][8] , \theRegs/managementDataOut[4][7] ,
         \theRegs/managementDataOut[4][6] , \theRegs/managementDataOut[4][5] ,
         \theRegs/managementDataOut[4][4] , \theRegs/managementDataOut[4][3] ,
         \theRegs/managementDataOut[4][2] , \theRegs/managementDataOut[4][1] ,
         \theRegs/managementDataOut[4][0] , \theRegs/managementDataOut[3][8] ,
         \theRegs/managementDataOut[3][7] , \theRegs/managementDataOut[3][6] ,
         \theRegs/managementDataOut[3][5] , \theRegs/managementDataOut[3][4] ,
         \theRegs/managementDataOut[3][3] , \theRegs/managementDataOut[3][2] ,
         \theRegs/managementDataOut[3][1] , \theRegs/managementDataOut[3][0] ,
         \theRegs/managementDataOut[2][8] , \theRegs/managementDataOut[2][7] ,
         \theRegs/managementDataOut[2][6] , \theRegs/managementDataOut[2][5] ,
         \theRegs/managementDataOut[2][4] , \theRegs/managementDataOut[2][3] ,
         \theRegs/managementDataOut[2][2] , \theRegs/managementDataOut[2][1] ,
         \theRegs/managementDataOut[2][0] , \theRegs/managementDataOut[1][8] ,
         \theRegs/managementDataOut[1][7] , \theRegs/managementDataOut[1][6] ,
         \theRegs/managementDataOut[1][5] , \theRegs/managementDataOut[1][4] ,
         \theRegs/managementDataOut[1][3] , \theRegs/managementDataOut[1][2] ,
         \theRegs/managementDataOut[1][1] , \theRegs/managementDataOut[1][0] ,
         \theRegs/managementDataOut[0][8] , \theRegs/managementDataOut[0][7] ,
         \theRegs/managementDataOut[0][6] , \theRegs/managementDataOut[0][5] ,
         \theRegs/managementDataOut[0][4] , \theRegs/managementDataOut[0][3] ,
         \theRegs/managementDataOut[0][2] , \theRegs/managementDataOut[0][1] ,
         \theRegs/managementDataOut[0][0] ,
         \theRegs/eachManagementReg[0].managementReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[0].managementReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[0].managementReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[0].managementReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[0].managementReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[0].managementReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[0].managementReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[0].managementReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[0].managementReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[1].managementReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[1].managementReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[1].managementReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[1].managementReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[1].managementReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[1].managementReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[1].managementReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[1].managementReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[1].managementReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[2].managementReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[2].managementReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[2].managementReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[2].managementReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[2].managementReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[2].managementReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[2].managementReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[2].managementReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[2].managementReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[3].managementReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[3].managementReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[3].managementReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[3].managementReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[3].managementReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[3].managementReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[3].managementReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[3].managementReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[3].managementReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[4].managementReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[4].managementReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[4].managementReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[4].managementReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[4].managementReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[4].managementReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[4].managementReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[4].managementReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[4].managementReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[5].managementReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[5].managementReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[5].managementReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[5].managementReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[5].managementReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[5].managementReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[5].managementReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[5].managementReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[5].managementReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[6].managementReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[6].managementReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[6].managementReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[6].managementReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[6].managementReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[6].managementReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[6].managementReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[6].managementReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[6].managementReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[7].managementReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[7].managementReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[7].managementReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[7].managementReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[7].managementReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[7].managementReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[7].managementReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[7].managementReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachManagementReg[7].managementReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[9].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[10].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[11].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[12].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[13].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[14].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[15].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[16].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[17].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[18].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[19].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[20].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[21].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[22].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[23].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[24].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[25].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[26].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[27].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[28].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[29].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[30].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[31].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[32].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[33].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[34].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[35].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[36].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[37].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[38].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[39].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[40].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[41].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[42].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[43].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[44].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[45].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[46].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[47].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[48].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[49].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[50].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[51].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[52].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[53].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[54].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[55].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[56].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[57].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[58].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[59].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[60].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[61].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[62].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[63].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[64].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[65].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[66].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[67].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[68].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[0].completionReg/eachEnDff[69].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[9].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[10].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[11].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[12].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[13].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[14].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[15].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[16].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[17].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[18].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[19].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[20].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[21].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[22].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[23].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[24].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[25].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[26].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[27].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[28].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[29].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[30].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[31].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[32].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[33].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[34].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[35].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[36].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[37].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[38].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[39].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[40].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[41].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[42].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[43].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[44].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[45].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[46].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[47].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[48].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[49].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[50].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[51].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[52].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[53].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[54].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[55].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[56].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[57].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[58].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[59].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[60].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[61].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[62].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[63].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[64].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[65].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[66].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[67].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[68].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[1].completionReg/eachEnDff[69].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[9].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[10].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[11].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[12].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[13].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[14].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[15].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[16].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[17].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[18].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[19].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[20].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[21].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[22].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[23].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[24].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[25].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[26].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[27].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[28].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[29].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[30].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[31].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[32].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[33].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[34].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[35].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[36].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[37].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[38].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[39].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[40].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[41].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[42].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[43].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[44].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[45].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[46].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[47].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[48].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[49].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[50].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[51].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[52].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[53].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[54].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[55].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[56].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[57].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[58].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[59].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[60].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[61].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[62].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[63].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[64].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[65].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[66].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[67].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[68].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[2].completionReg/eachEnDff[69].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[9].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[10].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[11].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[12].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[13].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[14].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[15].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[16].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[17].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[18].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[19].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[20].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[21].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[22].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[23].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[24].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[25].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[26].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[27].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[28].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[29].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[30].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[31].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[32].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[33].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[34].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[35].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[36].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[37].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[38].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[39].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[40].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[41].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[42].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[43].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[44].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[45].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[46].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[47].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[48].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[49].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[50].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[51].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[52].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[53].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[54].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[55].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[56].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[57].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[58].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[59].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[60].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[61].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[62].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[63].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[64].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[65].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[66].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[67].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[68].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[3].completionReg/eachEnDff[69].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[9].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[10].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[11].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[12].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[13].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[14].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[15].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[16].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[17].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[18].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[19].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[20].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[21].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[22].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[23].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[24].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[25].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[26].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[27].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[28].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[29].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[30].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[31].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[32].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[33].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[34].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[35].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[36].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[37].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[38].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[39].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[40].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[41].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[42].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[43].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[44].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[45].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[46].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[47].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[48].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[49].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[50].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[51].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[52].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[53].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[54].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[55].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[56].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[57].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[58].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[59].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[60].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[61].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[62].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[63].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[64].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[65].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[66].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[67].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[68].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[4].completionReg/eachEnDff[69].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[9].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[10].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[11].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[12].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[13].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[14].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[15].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[16].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[17].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[18].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[19].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[20].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[21].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[22].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[23].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[24].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[25].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[26].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[27].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[28].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[29].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[30].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[31].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[32].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[33].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[34].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[35].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[36].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[37].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[38].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[39].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[40].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[41].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[42].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[43].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[44].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[45].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[46].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[47].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[48].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[49].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[50].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[51].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[52].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[53].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[54].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[55].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[56].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[57].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[58].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[59].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[60].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[61].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[62].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[63].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[64].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[65].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[66].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[67].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[68].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[5].completionReg/eachEnDff[69].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[9].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[10].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[11].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[12].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[13].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[14].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[15].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[16].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[17].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[18].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[19].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[20].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[21].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[22].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[23].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[24].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[25].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[26].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[27].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[28].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[29].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[30].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[31].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[32].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[33].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[34].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[35].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[36].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[37].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[38].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[39].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[40].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[41].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[42].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[43].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[44].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[45].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[46].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[47].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[48].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[49].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[50].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[51].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[52].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[53].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[54].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[55].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[56].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[57].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[58].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[59].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[60].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[61].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[62].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[63].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[64].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[65].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[66].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[67].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[68].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[6].completionReg/eachEnDff[69].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[0].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[1].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[2].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[3].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[4].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[5].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[6].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[7].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[8].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[9].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[10].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[11].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[12].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[13].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[14].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[15].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[16].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[17].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[18].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[19].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[20].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[21].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[22].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[23].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[24].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[25].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[26].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[27].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[28].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[29].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[30].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[31].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[32].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[33].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[34].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[35].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[36].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[37].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[38].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[39].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[40].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[41].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[42].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[43].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[44].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[45].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[46].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[47].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[48].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[49].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[50].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[51].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[52].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[53].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[54].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[55].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[56].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[57].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[58].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[59].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[60].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[61].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[62].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[63].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[64].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[65].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[66].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[67].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[68].enDff/theFlop/N3 ,
         \theRegs/eachCompletionReg[7].completionReg/eachEnDff[69].enDff/theFlop/N3 ,
         \add_x_7/n1 , \add_x_6/n1 , n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2200, n2201, n2202, n2203, n2204, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2243, n2244, n2245, n2246, n2247, n2248, n2250,
         n2251, n2252, n2253, n2256, n2257, n2260, n2262, n2263, n2264, n2265,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2596, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117;
  wire   [2:0] tail;
  wire   [2:0] head;
  assign nextTail_o[3] = \add_x_6/n1 ;

  DFQD1 \headTailManager/headReset_reg  ( .D(n1407), .CP(clk_i), .Q(
        \headTailManager/headReset ) );
  DFQD1 \headTailManager/tail_reg[2]  ( .D(n1400), .CP(clk_i), .Q(tail[2]) );
  DFQD1 \theRegs/eachManagementReg[0].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[0][0] ) );
  DFQD1 \theRegs/eachManagementReg[0].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[0][1] ) );
  DFQD1 \theRegs/eachManagementReg[0].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[0][2] ) );
  DFQD1 \theRegs/eachManagementReg[0].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[0][3] ) );
  DFQD1 \theRegs/eachManagementReg[0].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[0][4] ) );
  DFQD1 \theRegs/eachManagementReg[0].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[0][5] ) );
  DFQD1 \theRegs/eachManagementReg[0].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[0][6] ) );
  DFQD1 \theRegs/eachManagementReg[0].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[0][7] ) );
  DFQD1 \theRegs/eachManagementReg[0].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[0][8] ) );
  DFQD1 \theRegs/eachManagementReg[1].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[1][0] ) );
  DFQD1 \theRegs/eachManagementReg[1].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[1][2] ) );
  DFQD1 \theRegs/eachManagementReg[1].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[1][3] ) );
  DFQD1 \theRegs/eachManagementReg[1].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[1][6] ) );
  DFQD1 \theRegs/eachManagementReg[1].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[1][8] ) );
  DFQD1 \theRegs/eachManagementReg[2].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[2][0] ) );
  DFQD1 \theRegs/eachManagementReg[2].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[2][1] ) );
  DFQD1 \theRegs/eachManagementReg[2].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[2][2] ) );
  DFQD1 \theRegs/eachManagementReg[2].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[2][3] ) );
  DFQD1 \theRegs/eachManagementReg[2].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[2][4] ) );
  DFQD1 \theRegs/eachManagementReg[2].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[2][5] ) );
  DFQD1 \theRegs/eachManagementReg[2].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[2][6] ) );
  DFQD1 \theRegs/eachManagementReg[2].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[2][7] ) );
  DFQD1 \theRegs/eachManagementReg[3].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[3][0] ) );
  DFQD1 \theRegs/eachManagementReg[3].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[3][1] ) );
  DFQD1 \theRegs/eachManagementReg[3].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[3][2] ) );
  DFQD1 \theRegs/eachManagementReg[3].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[3][3] ) );
  DFQD1 \theRegs/eachManagementReg[3].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[3][4] ) );
  DFQD1 \theRegs/eachManagementReg[3].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[3][5] ) );
  DFQD1 \theRegs/eachManagementReg[3].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[3][6] ) );
  DFQD1 \theRegs/eachManagementReg[3].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[3][7] ) );
  DFQD1 \theRegs/eachManagementReg[3].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[3][8] ) );
  DFQD1 \theRegs/eachManagementReg[4].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[4][0] ) );
  DFQD1 \theRegs/eachManagementReg[4].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[4][1] ) );
  DFQD1 \theRegs/eachManagementReg[4].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[4][2] ) );
  DFQD1 \theRegs/eachManagementReg[4].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[4][3] ) );
  DFQD1 \theRegs/eachManagementReg[4].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[4][4] ) );
  DFQD1 \theRegs/eachManagementReg[4].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[4][6] ) );
  DFQD1 \theRegs/eachManagementReg[5].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[5][0] ) );
  DFQD1 \theRegs/eachManagementReg[5].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[5][1] ) );
  DFQD1 \theRegs/eachManagementReg[5].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[5][2] ) );
  DFQD1 \theRegs/eachManagementReg[5].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[5][4] ) );
  DFQD1 \theRegs/eachManagementReg[5].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[5][5] ) );
  DFQD1 \theRegs/eachManagementReg[5].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[5][6] ) );
  DFQD1 \theRegs/eachManagementReg[5].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[5][7] ) );
  DFQD1 \theRegs/eachManagementReg[5].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[5][8] ) );
  DFQD1 \theRegs/eachManagementReg[6].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[6][0] ) );
  DFQD1 \theRegs/eachManagementReg[6].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[6][1] ) );
  DFQD1 \theRegs/eachManagementReg[6].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[6][2] ) );
  DFQD1 \theRegs/eachManagementReg[6].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[6][3] ) );
  DFQD1 \theRegs/eachManagementReg[6].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[6][4] ) );
  DFQD1 \theRegs/eachManagementReg[6].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[6][5] ) );
  DFQD1 \theRegs/eachManagementReg[6].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[6][6] ) );
  DFQD1 \theRegs/eachManagementReg[6].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[6][7] ) );
  DFQD1 \theRegs/eachManagementReg[6].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[6][8] ) );
  DFQD1 \theRegs/eachManagementReg[7].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[7][1] ) );
  DFQD1 \theRegs/eachManagementReg[7].managementReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[7][2] ) );
  DFQD1 \theRegs/eachManagementReg[7].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[7][3] ) );
  DFQD1 \theRegs/eachManagementReg[7].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[7][4] ) );
  DFQD1 \theRegs/eachManagementReg[7].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[7][5] ) );
  DFQD1 \theRegs/eachManagementReg[7].managementReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[7][6] ) );
  DFQD1 \theRegs/eachManagementReg[7].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[7][7] ) );
  DFQD1 \theRegs/eachManagementReg[7].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[7][8] ) );
  DFQD1 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[65].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][65] ) );
  DFQD1 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[66].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][66] ) );
  DFQD1 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[67].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][67] ) );
  DFQD1 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[68].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][68] ) );
  DFQD1 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[69].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][69] ) );
  DFQD1 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[65].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][65] ) );
  DFQD1 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[66].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][66] ) );
  DFQD1 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[67].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][67] ) );
  DFQD1 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[68].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][68] ) );
  DFQD1 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[69].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][69] ) );
  DFQD1 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[65].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][65] ) );
  DFQD1 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[66].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][66] ) );
  DFQD1 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[67].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][67] ) );
  DFQD1 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[68].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][68] ) );
  DFQD1 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[69].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][69] ) );
  DFQD1 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[65].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][65] ) );
  DFQD1 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[66].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][66] ) );
  DFQD1 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[67].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][67] ) );
  DFQD1 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[68].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][68] ) );
  DFQD1 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[69].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][69] ) );
  DFQD1 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[65].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][65] ) );
  DFQD1 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[66].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][66] ) );
  DFQD1 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[67].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][67] ) );
  DFQD1 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[68].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][68] ) );
  DFQD1 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[69].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][69] ) );
  DFQD1 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[65].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][65] ) );
  DFQD1 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[66].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][66] ) );
  DFQD1 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[67].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][67] ) );
  DFQD1 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[68].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][68] ) );
  DFQD1 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[69].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][69] ) );
  DFQD1 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[65].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][65] ) );
  DFQD1 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[66].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][66] ) );
  DFQD1 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[67].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][67] ) );
  DFQD1 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[68].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][68] ) );
  DFQD1 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[69].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][69] ) );
  DFQD1 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[65].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[65].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][65] ) );
  DFQD1 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[66].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[66].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][66] ) );
  DFQD1 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[67].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[67].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][67] ) );
  DFQD1 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[68].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[68].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][68] ) );
  DFQD1 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[69].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[69].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][69] ) );
  ND2D0 U2314 ( .A1(n3229), .A2(n3225), .ZN(n2871) );
  AO22D0 U2333 ( .A1(n3210), .A2(n3677), .B1(
        \theRegs/completionDataOut[0][69] ), .B2(n3520), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[69].enDff/theFlop/N3 ) );
  AO22D0 U2334 ( .A1(n3209), .A2(n3711), .B1(n3648), .B2(
        \theRegs/completionDataOut[0][68] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[68].enDff/theFlop/N3 ) );
  AO22D0 U2335 ( .A1(n3208), .A2(n3677), .B1(n3468), .B2(
        \theRegs/completionDataOut[0][67] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[67].enDff/theFlop/N3 ) );
  AO22D0 U2336 ( .A1(n3207), .A2(n3559), .B1(n3468), .B2(
        \theRegs/completionDataOut[0][66] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[66].enDff/theFlop/N3 ) );
  AO22D0 U2337 ( .A1(n3198), .A2(n3663), .B1(n3622), .B2(
        \theRegs/completionDataOut[0][57] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[57].enDff/theFlop/N3 ) );
  AO22D0 U2338 ( .A1(n4050), .A2(n3711), .B1(n3766), .B2(
        \theRegs/completionDataOut[0][59] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[59].enDff/theFlop/N3 ) );
  AO22D0 U2339 ( .A1(n4052), .A2(n3845), .B1(n3796), .B2(
        \theRegs/completionDataOut[0][58] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[58].enDff/theFlop/N3 ) );
  AO22D0 U2340 ( .A1(n4073), .A2(n3586), .B1(n3628), .B2(
        \theRegs/completionDataOut[0][61] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[61].enDff/theFlop/N3 ) );
  AO22D0 U2341 ( .A1(n3204), .A2(n3677), .B1(n3468), .B2(
        \theRegs/completionDataOut[0][63] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[63].enDff/theFlop/N3 ) );
  AO22D0 U2342 ( .A1(n3203), .A2(n3475), .B1(n3448), .B2(
        \theRegs/completionDataOut[0][62] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[62].enDff/theFlop/N3 ) );
  AO22D0 U2343 ( .A1(n3205), .A2(n3677), .B1(n3628), .B2(
        \theRegs/completionDataOut[0][64] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[64].enDff/theFlop/N3 ) );
  AO22D0 U2344 ( .A1(n3201), .A2(n3475), .B1(n3448), .B2(
        \theRegs/completionDataOut[0][60] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[60].enDff/theFlop/N3 ) );
  AO22D0 U2345 ( .A1(n4082), .A2(n3803), .B1(n3864), .B2(
        \theRegs/completionDataOut[0][56] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[56].enDff/theFlop/N3 ) );
  AO22D0 U2346 ( .A1(n4074), .A2(n3921), .B1(n3622), .B2(
        \theRegs/completionDataOut[0][55] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[55].enDff/theFlop/N3 ) );
  AO22D0 U2347 ( .A1(n3195), .A2(n4020), .B1(n3757), .B2(
        \theRegs/completionDataOut[0][54] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[54].enDff/theFlop/N3 ) );
  AO22D0 U2348 ( .A1(n3206), .A2(n3812), .B1(n3766), .B2(
        \theRegs/completionDataOut[0][65] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[65].enDff/theFlop/N3 ) );
  AO22D0 U2350 ( .A1(n3180), .A2(n3559), .B1(n3520), .B2(
        \theRegs/completionDataOut[0][39] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[39].enDff/theFlop/N3 ) );
  AO22D0 U2351 ( .A1(n4107), .A2(n4020), .B1(n4003), .B2(
        \theRegs/completionDataOut[0][47] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[47].enDff/theFlop/N3 ) );
  AO22D0 U2352 ( .A1(n3163), .A2(n3663), .B1(n3727), .B2(
        \theRegs/completionDataOut[0][22] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[22].enDff/theFlop/N3 ) );
  AO22D0 U2353 ( .A1(n3186), .A2(n3559), .B1(n3468), .B2(
        \theRegs/completionDataOut[0][45] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[45].enDff/theFlop/N3 ) );
  AO22D0 U2354 ( .A1(n3185), .A2(n3475), .B1(n3448), .B2(
        \theRegs/completionDataOut[0][44] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[44].enDff/theFlop/N3 ) );
  AO22D0 U2355 ( .A1(n4100), .A2(n3845), .B1(n3907), .B2(
        \theRegs/completionDataOut[0][43] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[43].enDff/theFlop/N3 ) );
  AO22D0 U2356 ( .A1(n4095), .A2(n3812), .B1(n3541), .B2(
        \theRegs/completionDataOut[0][42] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[42].enDff/theFlop/N3 ) );
  AO22D0 U2357 ( .A1(n4097), .A2(n3586), .B1(n3541), .B2(
        \theRegs/completionDataOut[0][41] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[41].enDff/theFlop/N3 ) );
  AO22D0 U2358 ( .A1(n4101), .A2(n3845), .B1(n3796), .B2(
        \theRegs/completionDataOut[0][40] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[40].enDff/theFlop/N3 ) );
  AO22D0 U2359 ( .A1(n4102), .A2(n3956), .B1(n3893), .B2(
        \theRegs/completionDataOut[0][49] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[49].enDff/theFlop/N3 ) );
  AO22D0 U2360 ( .A1(n3189), .A2(n3803), .B1(n3757), .B2(
        \theRegs/completionDataOut[0][48] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[48].enDff/theFlop/N3 ) );
  AO22D0 U2361 ( .A1(n4067), .A2(n3956), .B1(n3893), .B2(
        \theRegs/completionDataOut[0][52] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[52].enDff/theFlop/N3 ) );
  AO22D0 U2362 ( .A1(n4076), .A2(n3956), .B1(n3893), .B2(
        \theRegs/completionDataOut[0][46] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[46].enDff/theFlop/N3 ) );
  AO22D0 U2363 ( .A1(n3191), .A2(n3803), .B1(n3757), .B2(
        \theRegs/completionDataOut[0][50] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[50].enDff/theFlop/N3 ) );
  AO22D0 U2364 ( .A1(n4091), .A2(n3812), .B1(n3541), .B2(
        \theRegs/completionDataOut[0][10] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[10].enDff/theFlop/N3 ) );
  AO22D0 U2365 ( .A1(n3150), .A2(n3812), .B1(n3766), .B2(
        \theRegs/completionDataOut[0][9] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[9].enDff/theFlop/N3 ) );
  AO22D0 U2366 ( .A1(n3149), .A2(n3711), .B1(n3648), .B2(
        \theRegs/completionDataOut[0][8] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U2367 ( .A1(n3148), .A2(n3475), .B1(n3309), .B2(
        \theRegs/completionDataOut[0][7] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U2368 ( .A1(n3147), .A2(n3559), .B1(n3468), .B2(
        \theRegs/completionDataOut[0][6] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U2369 ( .A1(n3146), .A2(n3475), .B1(n3448), .B2(
        \theRegs/completionDataOut[0][5] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U2370 ( .A1(n3145), .A2(n3559), .B1(n3520), .B2(
        \theRegs/completionDataOut[0][4] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U2371 ( .A1(n3144), .A2(n3586), .B1(n3541), .B2(
        \theRegs/completionDataOut[0][3] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U2372 ( .A1(n3143), .A2(n3711), .B1(n3648), .B2(
        \theRegs/completionDataOut[0][2] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U2373 ( .A1(n3142), .A2(n3586), .B1(n3628), .B2(
        \theRegs/completionDataOut[0][1] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U2374 ( .A1(n4075), .A2(n3845), .B1(n3796), .B2(
        \theRegs/completionDataOut[0][0] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U2375 ( .A1(n4063), .A2(n3845), .B1(n3796), .B2(
        \theRegs/completionDataOut[0][38] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[38].enDff/theFlop/N3 ) );
  AO22D0 U2376 ( .A1(n4077), .A2(n3812), .B1(n3541), .B2(
        \theRegs/completionDataOut[0][37] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[37].enDff/theFlop/N3 ) );
  AO22D0 U2377 ( .A1(n4072), .A2(n3960), .B1(n3907), .B2(
        \theRegs/completionDataOut[0][36] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[36].enDff/theFlop/N3 ) );
  AO22D0 U2378 ( .A1(n4106), .A2(n3960), .B1(n3907), .B2(
        \theRegs/completionDataOut[0][35] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[35].enDff/theFlop/N3 ) );
  AO22D0 U2379 ( .A1(n3192), .A2(n3663), .B1(n3727), .B2(
        \theRegs/completionDataOut[0][51] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[51].enDff/theFlop/N3 ) );
  AO22D0 U2380 ( .A1(n4045), .A2(n3586), .B1(n3541), .B2(
        \theRegs/completionDataOut[0][33] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[33].enDff/theFlop/N3 ) );
  AO22D0 U2381 ( .A1(n3173), .A2(n3559), .B1(n3520), .B2(
        \theRegs/completionDataOut[0][32] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[32].enDff/theFlop/N3 ) );
  AO22D0 U2382 ( .A1(n4047), .A2(n4020), .B1(n3757), .B2(
        \theRegs/completionDataOut[0][31] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[31].enDff/theFlop/N3 ) );
  AO22D0 U2383 ( .A1(n4051), .A2(n3956), .B1(n3893), .B2(
        \theRegs/completionDataOut[0][30] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[30].enDff/theFlop/N3 ) );
  AO22D0 U2384 ( .A1(n4105), .A2(n3781), .B1(n3588), .B2(
        \theRegs/completionDataOut[0][29] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[29].enDff/theFlop/N3 ) );
  AO22D0 U2385 ( .A1(n4103), .A2(n3956), .B1(n3893), .B2(
        \theRegs/completionDataOut[0][28] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[28].enDff/theFlop/N3 ) );
  AO22D0 U2386 ( .A1(n4109), .A2(n3803), .B1(n3864), .B2(
        \theRegs/completionDataOut[0][27] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[27].enDff/theFlop/N3 ) );
  AO22D0 U2387 ( .A1(n4110), .A2(n3663), .B1(n3622), .B2(
        \theRegs/completionDataOut[0][26] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[26].enDff/theFlop/N3 ) );
  AO22D0 U2388 ( .A1(n4111), .A2(n4020), .B1(n3757), .B2(
        \theRegs/completionDataOut[0][25] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[25].enDff/theFlop/N3 ) );
  AO22D0 U2389 ( .A1(n4098), .A2(n3803), .B1(n3757), .B2(
        \theRegs/completionDataOut[0][24] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[24].enDff/theFlop/N3 ) );
  AO22D0 U2390 ( .A1(n3164), .A2(n3803), .B1(n3864), .B2(
        \theRegs/completionDataOut[0][23] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[23].enDff/theFlop/N3 ) );
  AO22D0 U2391 ( .A1(n3194), .A2(n3310), .B1(n3308), .B2(
        \theRegs/completionDataOut[0][53] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[53].enDff/theFlop/N3 ) );
  AO22D0 U2394 ( .A1(n3162), .A2(n3310), .B1(n3308), .B2(
        \theRegs/completionDataOut[0][21] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[21].enDff/theFlop/N3 ) );
  AO22D0 U2395 ( .A1(n3161), .A2(n3781), .B1(n3588), .B2(
        \theRegs/completionDataOut[0][20] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[20].enDff/theFlop/N3 ) );
  AO22D0 U2396 ( .A1(n4044), .A2(n3663), .B1(n3727), .B2(
        \theRegs/completionDataOut[0][19] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[19].enDff/theFlop/N3 ) );
  AO22D0 U2397 ( .A1(n4114), .A2(n3921), .B1(n3622), .B2(
        \theRegs/completionDataOut[0][18] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[18].enDff/theFlop/N3 ) );
  AO22D0 U2398 ( .A1(n3175), .A2(n3711), .B1(n3648), .B2(
        \theRegs/completionDataOut[0][34] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[34].enDff/theFlop/N3 ) );
  AO22D0 U2401 ( .A1(n3157), .A2(n3781), .B1(n3588), .B2(
        \theRegs/completionDataOut[0][16] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[16].enDff/theFlop/N3 ) );
  AO22D0 U2402 ( .A1(n4053), .A2(n3921), .B1(n3622), .B2(
        \theRegs/completionDataOut[0][15] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[15].enDff/theFlop/N3 ) );
  AO22D0 U2403 ( .A1(n3155), .A2(n3310), .B1(n3588), .B2(
        \theRegs/completionDataOut[0][14] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[14].enDff/theFlop/N3 ) );
  AO22D0 U2404 ( .A1(n4055), .A2(n3663), .B1(n3622), .B2(
        \theRegs/completionDataOut[0][13] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[13].enDff/theFlop/N3 ) );
  AO22D0 U2405 ( .A1(n4056), .A2(n3956), .B1(n3893), .B2(
        \theRegs/completionDataOut[0][12] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[12].enDff/theFlop/N3 ) );
  AO22D0 U2406 ( .A1(n3152), .A2(n3475), .B1(n3448), .B2(
        \theRegs/completionDataOut[0][11] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[11].enDff/theFlop/N3 ) );
  AO22D0 U2408 ( .A1(n3158), .A2(n3781), .B1(n3588), .B2(
        \theRegs/completionDataOut[0][17] ), .Z(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[17].enDff/theFlop/N3 ) );
  AO22D0 U2417 ( .A1(n3210), .A2(n3450), .B1(
        \theRegs/completionDataOut[4][69] ), .B2(n3780), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[69].enDff/theFlop/N3 ) );
  AO22D0 U2418 ( .A1(n4069), .A2(n3460), .B1(n3849), .B2(
        \theRegs/completionDataOut[4][67] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[67].enDff/theFlop/N3 ) );
  AO22D0 U2419 ( .A1(n4060), .A2(n3401), .B1(n3780), .B2(
        \theRegs/completionDataOut[4][66] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[66].enDff/theFlop/N3 ) );
  AO22D0 U2420 ( .A1(n3209), .A2(n3387), .B1(n3713), .B2(
        \theRegs/completionDataOut[4][68] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[68].enDff/theFlop/N3 ) );
  AO22D0 U2421 ( .A1(n3196), .A2(n3871), .B1(n3925), .B2(
        \theRegs/completionDataOut[4][55] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[55].enDff/theFlop/N3 ) );
  AO22D0 U2422 ( .A1(n3205), .A2(n3512), .B1(n3853), .B2(
        \theRegs/completionDataOut[4][64] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[64].enDff/theFlop/N3 ) );
  AO22D0 U2423 ( .A1(n3204), .A2(n3512), .B1(n3853), .B2(
        \theRegs/completionDataOut[4][63] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[63].enDff/theFlop/N3 ) );
  AO22D0 U2424 ( .A1(n4064), .A2(n3589), .B1(n3849), .B2(
        \theRegs/completionDataOut[4][65] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[65].enDff/theFlop/N3 ) );
  AO22D0 U2425 ( .A1(n4073), .A2(n3401), .B1(n3825), .B2(
        \theRegs/completionDataOut[4][61] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[61].enDff/theFlop/N3 ) );
  AO22D0 U2426 ( .A1(n3201), .A2(n3387), .B1(n3780), .B2(
        \theRegs/completionDataOut[4][60] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[60].enDff/theFlop/N3 ) );
  AO22D0 U2427 ( .A1(n4050), .A2(n3460), .B1(n3849), .B2(
        \theRegs/completionDataOut[4][59] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[59].enDff/theFlop/N3 ) );
  AO22D0 U2428 ( .A1(n4052), .A2(n3460), .B1(n3849), .B2(
        \theRegs/completionDataOut[4][58] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[58].enDff/theFlop/N3 ) );
  AO22D0 U2429 ( .A1(n4086), .A2(n3955), .B1(n4015), .B2(
        \theRegs/completionDataOut[4][57] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[57].enDff/theFlop/N3 ) );
  AO22D0 U2430 ( .A1(n3197), .A2(n3612), .B1(n3657), .B2(
        \theRegs/completionDataOut[4][56] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[56].enDff/theFlop/N3 ) );
  AO22D0 U2431 ( .A1(n3203), .A2(n3589), .B1(n3849), .B2(
        \theRegs/completionDataOut[4][62] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[62].enDff/theFlop/N3 ) );
  AO22D0 U2432 ( .A1(n3195), .A2(n3612), .B1(n3657), .B2(
        \theRegs/completionDataOut[4][54] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[54].enDff/theFlop/N3 ) );
  AO22D0 U2434 ( .A1(n4075), .A2(n3589), .B1(n3969), .B2(
        \theRegs/completionDataOut[4][0] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U2435 ( .A1(n3194), .A2(n3612), .B1(n3657), .B2(
        \theRegs/completionDataOut[4][53] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[53].enDff/theFlop/N3 ) );
  AO22D0 U2436 ( .A1(n3193), .A2(n3871), .B1(n3925), .B2(
        \theRegs/completionDataOut[4][52] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[52].enDff/theFlop/N3 ) );
  AO22D0 U2438 ( .A1(n3192), .A2(n3612), .B1(n3657), .B2(
        \theRegs/completionDataOut[4][51] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[51].enDff/theFlop/N3 ) );
  AO22D0 U2439 ( .A1(n3191), .A2(n3760), .B1(n3806), .B2(
        \theRegs/completionDataOut[4][50] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[50].enDff/theFlop/N3 ) );
  AO22D0 U2440 ( .A1(n3190), .A2(n4000), .B1(n4037), .B2(
        \theRegs/completionDataOut[4][49] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[49].enDff/theFlop/N3 ) );
  AO22D0 U2441 ( .A1(n3189), .A2(n3760), .B1(n3806), .B2(
        \theRegs/completionDataOut[4][48] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[48].enDff/theFlop/N3 ) );
  AO22D0 U2442 ( .A1(n4107), .A2(n3955), .B1(n4015), .B2(
        \theRegs/completionDataOut[4][47] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[47].enDff/theFlop/N3 ) );
  AO22D0 U2443 ( .A1(n3187), .A2(n3732), .B1(n3787), .B2(
        \theRegs/completionDataOut[4][46] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[46].enDff/theFlop/N3 ) );
  AO22D0 U2444 ( .A1(n4094), .A2(n3401), .B1(n3780), .B2(
        \theRegs/completionDataOut[4][45] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[45].enDff/theFlop/N3 ) );
  AO22D0 U2445 ( .A1(n4108), .A2(n3426), .B1(n3914), .B2(
        \theRegs/completionDataOut[4][44] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[44].enDff/theFlop/N3 ) );
  AO22D0 U2446 ( .A1(n4100), .A2(n3387), .B1(n3713), .B2(
        \theRegs/completionDataOut[4][43] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[43].enDff/theFlop/N3 ) );
  AO22D0 U2447 ( .A1(n4095), .A2(n3401), .B1(n3780), .B2(
        \theRegs/completionDataOut[4][42] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[42].enDff/theFlop/N3 ) );
  AO22D0 U2448 ( .A1(n4097), .A2(n3401), .B1(n3780), .B2(
        \theRegs/completionDataOut[4][41] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[41].enDff/theFlop/N3 ) );
  AO22D0 U2449 ( .A1(n3181), .A2(n3426), .B1(n3914), .B2(
        \theRegs/completionDataOut[4][40] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[40].enDff/theFlop/N3 ) );
  AO22D0 U2450 ( .A1(n4081), .A2(n3426), .B1(n3914), .B2(
        \theRegs/completionDataOut[4][39] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[39].enDff/theFlop/N3 ) );
  AO22D0 U2451 ( .A1(n3179), .A2(n3426), .B1(n3914), .B2(
        \theRegs/completionDataOut[4][38] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[38].enDff/theFlop/N3 ) );
  AO22D0 U2452 ( .A1(n4077), .A2(n3539), .B1(n3969), .B2(
        \theRegs/completionDataOut[4][37] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[37].enDff/theFlop/N3 ) );
  AO22D0 U2453 ( .A1(n3177), .A2(n3539), .B1(n3969), .B2(
        \theRegs/completionDataOut[4][36] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[36].enDff/theFlop/N3 ) );
  AO22D0 U2455 ( .A1(n4106), .A2(n3539), .B1(n3969), .B2(
        \theRegs/completionDataOut[4][35] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[35].enDff/theFlop/N3 ) );
  AO22D0 U2456 ( .A1(n4098), .A2(n3955), .B1(n4015), .B2(
        \theRegs/completionDataOut[4][24] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[24].enDff/theFlop/N3 ) );
  AO22D0 U2457 ( .A1(n4104), .A2(n3539), .B1(n3890), .B2(
        \theRegs/completionDataOut[4][34] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[34].enDff/theFlop/N3 ) );
  AO22D0 U2459 ( .A1(n3174), .A2(n3342), .B1(n3330), .B2(
        \theRegs/completionDataOut[4][33] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[33].enDff/theFlop/N3 ) );
  AO22D0 U2460 ( .A1(n4046), .A2(n3539), .B1(n3890), .B2(
        \theRegs/completionDataOut[4][32] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[32].enDff/theFlop/N3 ) );
  AO22D0 U2461 ( .A1(n4047), .A2(n3401), .B1(n3825), .B2(
        \theRegs/completionDataOut[4][31] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[31].enDff/theFlop/N3 ) );
  AO22D0 U2462 ( .A1(n4051), .A2(n3539), .B1(n3890), .B2(
        \theRegs/completionDataOut[4][30] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[30].enDff/theFlop/N3 ) );
  AO22D0 U2463 ( .A1(n4105), .A2(n3760), .B1(n3806), .B2(
        \theRegs/completionDataOut[4][29] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[29].enDff/theFlop/N3 ) );
  AO22D0 U2464 ( .A1(n4103), .A2(n3955), .B1(n4015), .B2(
        \theRegs/completionDataOut[4][28] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[28].enDff/theFlop/N3 ) );
  AO22D0 U2465 ( .A1(n4109), .A2(n4000), .B1(n4037), .B2(
        \theRegs/completionDataOut[4][27] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[27].enDff/theFlop/N3 ) );
  AO22D0 U2466 ( .A1(n4110), .A2(n3955), .B1(n4015), .B2(
        \theRegs/completionDataOut[4][26] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[26].enDff/theFlop/N3 ) );
  AO22D0 U2467 ( .A1(n4111), .A2(n3760), .B1(n3806), .B2(
        \theRegs/completionDataOut[4][25] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[25].enDff/theFlop/N3 ) );
  AO22D0 U2468 ( .A1(n4091), .A2(n3426), .B1(n3853), .B2(
        \theRegs/completionDataOut[4][10] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[10].enDff/theFlop/N3 ) );
  AO22D0 U2469 ( .A1(n3164), .A2(n3760), .B1(n3806), .B2(
        \theRegs/completionDataOut[4][23] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[23].enDff/theFlop/N3 ) );
  AO22D0 U2470 ( .A1(n3163), .A2(n3732), .B1(n3787), .B2(
        \theRegs/completionDataOut[4][22] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[22].enDff/theFlop/N3 ) );
  AO22D0 U2471 ( .A1(n4112), .A2(n3341), .B1(n3329), .B2(
        \theRegs/completionDataOut[4][21] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[21].enDff/theFlop/N3 ) );
  AO22D0 U2472 ( .A1(n4113), .A2(n3955), .B1(n4015), .B2(
        \theRegs/completionDataOut[4][20] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[20].enDff/theFlop/N3 ) );
  AO22D0 U2473 ( .A1(n4044), .A2(n3341), .B1(n3329), .B2(
        \theRegs/completionDataOut[4][19] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[19].enDff/theFlop/N3 ) );
  AO22D0 U2474 ( .A1(n3159), .A2(n3612), .B1(n3657), .B2(
        \theRegs/completionDataOut[4][18] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[18].enDff/theFlop/N3 ) );
  AO22D0 U2476 ( .A1(n4048), .A2(n4000), .B1(n4037), .B2(
        \theRegs/completionDataOut[4][17] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[17].enDff/theFlop/N3 ) );
  AO22D0 U2477 ( .A1(n4049), .A2(n3871), .B1(n3925), .B2(
        \theRegs/completionDataOut[4][16] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[16].enDff/theFlop/N3 ) );
  AO22D0 U2480 ( .A1(n3156), .A2(n3612), .B1(n3657), .B2(
        \theRegs/completionDataOut[4][15] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[15].enDff/theFlop/N3 ) );
  AO22D0 U2481 ( .A1(n3145), .A2(n3512), .B1(n3853), .B2(
        \theRegs/completionDataOut[4][4] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U2482 ( .A1(n3142), .A2(n3450), .B1(n3825), .B2(
        \theRegs/completionDataOut[4][1] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U2483 ( .A1(n3143), .A2(n3460), .B1(n3988), .B2(
        \theRegs/completionDataOut[4][2] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U2484 ( .A1(n4054), .A2(n4000), .B1(n4037), .B2(
        \theRegs/completionDataOut[4][14] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[14].enDff/theFlop/N3 ) );
  AO22D0 U2485 ( .A1(n4055), .A2(n3760), .B1(n3806), .B2(
        \theRegs/completionDataOut[4][13] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[13].enDff/theFlop/N3 ) );
  AO22D0 U2486 ( .A1(n4056), .A2(n3341), .B1(n3329), .B2(
        \theRegs/completionDataOut[4][12] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[12].enDff/theFlop/N3 ) );
  AO22D0 U2487 ( .A1(n3152), .A2(n3450), .B1(n3825), .B2(
        \theRegs/completionDataOut[4][11] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[11].enDff/theFlop/N3 ) );
  AO22D0 U2488 ( .A1(n3146), .A2(n3387), .B1(n3713), .B2(
        \theRegs/completionDataOut[4][5] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U2489 ( .A1(n3150), .A2(n3387), .B1(n3713), .B2(
        \theRegs/completionDataOut[4][9] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[9].enDff/theFlop/N3 ) );
  AO22D0 U2490 ( .A1(n3149), .A2(n3426), .B1(n3914), .B2(
        \theRegs/completionDataOut[4][8] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U2491 ( .A1(n4090), .A2(n3450), .B1(n3825), .B2(
        \theRegs/completionDataOut[4][7] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U2492 ( .A1(n3147), .A2(n3387), .B1(n3713), .B2(
        \theRegs/completionDataOut[4][6] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U2493 ( .A1(n3144), .A2(n3450), .B1(n3825), .B2(
        \theRegs/completionDataOut[4][3] ), .Z(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U2501 ( .A1(n4068), .A2(n3994), .B1(
        \theRegs/completionDataOut[2][69] ), .B2(n3364), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[69].enDff/theFlop/N3 ) );
  AO22D0 U2502 ( .A1(n4059), .A2(n3897), .B1(n3388), .B2(
        \theRegs/completionDataOut[2][68] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[68].enDff/theFlop/N3 ) );
  AO22D0 U2503 ( .A1(n4069), .A2(n3994), .B1(n3427), .B2(
        \theRegs/completionDataOut[2][67] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[67].enDff/theFlop/N3 ) );
  AO22D0 U2504 ( .A1(n4060), .A2(n3701), .B1(n3361), .B2(
        \theRegs/completionDataOut[2][66] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[66].enDff/theFlop/N3 ) );
  AO22D0 U2505 ( .A1(n3202), .A2(n3328), .B1(n3315), .B2(
        \theRegs/completionDataOut[6][61] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[61].enDff/theFlop/N3 ) );
  AO22D0 U2506 ( .A1(n3204), .A2(n3710), .B1(n3315), .B2(
        \theRegs/completionDataOut[6][63] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[63].enDff/theFlop/N3 ) );
  AO22D0 U2507 ( .A1(n4065), .A2(n3844), .B1(n3998), .B2(
        \theRegs/completionDataOut[6][62] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[62].enDff/theFlop/N3 ) );
  AO22D0 U2508 ( .A1(n4085), .A2(n4022), .B1(n3807), .B2(
        \theRegs/completionDataOut[6][54] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[54].enDff/theFlop/N3 ) );
  AO22D0 U2509 ( .A1(n3201), .A2(n3710), .B1(n3315), .B2(
        \theRegs/completionDataOut[6][60] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[60].enDff/theFlop/N3 ) );
  AO22D0 U2510 ( .A1(n3205), .A2(n3710), .B1(n3315), .B2(
        \theRegs/completionDataOut[6][64] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[64].enDff/theFlop/N3 ) );
  AO22D0 U2511 ( .A1(n3199), .A2(n3827), .B1(n3970), .B2(
        \theRegs/completionDataOut[6][58] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[58].enDff/theFlop/N3 ) );
  AO22D0 U2512 ( .A1(n4086), .A2(n4022), .B1(n3859), .B2(
        \theRegs/completionDataOut[6][57] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[57].enDff/theFlop/N3 ) );
  AO22D0 U2513 ( .A1(n3197), .A2(n3709), .B1(n3859), .B2(
        \theRegs/completionDataOut[6][56] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[56].enDff/theFlop/N3 ) );
  AO22D0 U2514 ( .A1(n4074), .A2(n3709), .B1(n3859), .B2(
        \theRegs/completionDataOut[6][55] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[55].enDff/theFlop/N3 ) );
  AO22D0 U2515 ( .A1(n4050), .A2(n3749), .B1(n4018), .B2(
        \theRegs/completionDataOut[6][59] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[59].enDff/theFlop/N3 ) );
  AO22D0 U2516 ( .A1(n3206), .A2(n3827), .B1(n3970), .B2(
        \theRegs/completionDataOut[6][65] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[65].enDff/theFlop/N3 ) );
  AO22D0 U2517 ( .A1(n3210), .A2(n3844), .B1(
        \theRegs/completionDataOut[6][69] ), .B2(n4018), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[69].enDff/theFlop/N3 ) );
  AO22D0 U2518 ( .A1(n4059), .A2(n3844), .B1(n3998), .B2(
        \theRegs/completionDataOut[6][68] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[68].enDff/theFlop/N3 ) );
  AO22D0 U2519 ( .A1(n4069), .A2(n3844), .B1(n3998), .B2(
        \theRegs/completionDataOut[6][67] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[67].enDff/theFlop/N3 ) );
  AO22D0 U2520 ( .A1(n4060), .A2(n3749), .B1(n3848), .B2(
        \theRegs/completionDataOut[6][66] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[66].enDff/theFlop/N3 ) );
  AO22D0 U2522 ( .A1(n3195), .A2(n3701), .B1(n3351), .B2(
        \theRegs/completionDataOut[2][54] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[54].enDff/theFlop/N3 ) );
  AO22D0 U2523 ( .A1(n4064), .A2(n3897), .B1(n3417), .B2(
        \theRegs/completionDataOut[2][65] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[65].enDff/theFlop/N3 ) );
  AO22D0 U2524 ( .A1(n3205), .A2(n3869), .B1(n3351), .B2(
        \theRegs/completionDataOut[2][64] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[64].enDff/theFlop/N3 ) );
  AO22D0 U2525 ( .A1(n3204), .A2(n3897), .B1(n3388), .B2(
        \theRegs/completionDataOut[2][63] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[63].enDff/theFlop/N3 ) );
  AO22D0 U2526 ( .A1(n3203), .A2(n3802), .B1(n3364), .B2(
        \theRegs/completionDataOut[2][62] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[62].enDff/theFlop/N3 ) );
  AO22D0 U2527 ( .A1(n3202), .A2(n3785), .B1(n3349), .B2(
        \theRegs/completionDataOut[2][61] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[61].enDff/theFlop/N3 ) );
  AO22D0 U2528 ( .A1(n3201), .A2(n3869), .B1(n3351), .B2(
        \theRegs/completionDataOut[2][60] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[60].enDff/theFlop/N3 ) );
  AO22D0 U2529 ( .A1(n3200), .A2(n3339), .B1(n3349), .B2(
        \theRegs/completionDataOut[2][59] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[59].enDff/theFlop/N3 ) );
  AO22D0 U2530 ( .A1(n4052), .A2(n3949), .B1(n3427), .B2(
        \theRegs/completionDataOut[2][58] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[58].enDff/theFlop/N3 ) );
  AO22D0 U2531 ( .A1(n3198), .A2(n3701), .B1(n3351), .B2(
        \theRegs/completionDataOut[2][57] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[57].enDff/theFlop/N3 ) );
  AO22D0 U2532 ( .A1(n3197), .A2(n3785), .B1(n3349), .B2(
        \theRegs/completionDataOut[2][56] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[56].enDff/theFlop/N3 ) );
  AO22D0 U2533 ( .A1(n3196), .A2(n3339), .B1(n3349), .B2(
        \theRegs/completionDataOut[2][55] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[55].enDff/theFlop/N3 ) );
  AO22D0 U2535 ( .A1(n4046), .A2(n3915), .B1(n3623), .B2(
        \theRegs/completionDataOut[6][32] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[32].enDff/theFlop/N3 ) );
  AO22D0 U2536 ( .A1(n3187), .A2(n3915), .B1(n3623), .B2(
        \theRegs/completionDataOut[6][46] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[46].enDff/theFlop/N3 ) );
  AO22D0 U2537 ( .A1(n4067), .A2(n4022), .B1(n3807), .B2(
        \theRegs/completionDataOut[6][52] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[52].enDff/theFlop/N3 ) );
  AO22D0 U2538 ( .A1(n4057), .A2(n3709), .B1(n3859), .B2(
        \theRegs/completionDataOut[6][51] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[51].enDff/theFlop/N3 ) );
  AO22D0 U2539 ( .A1(n4058), .A2(n4022), .B1(n3807), .B2(
        \theRegs/completionDataOut[6][50] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[50].enDff/theFlop/N3 ) );
  AO22D0 U2540 ( .A1(n3183), .A2(n3710), .B1(n3970), .B2(
        \theRegs/completionDataOut[6][42] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[42].enDff/theFlop/N3 ) );
  AO22D0 U2541 ( .A1(n4097), .A2(n3710), .B1(n3970), .B2(
        \theRegs/completionDataOut[6][41] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[41].enDff/theFlop/N3 ) );
  AO22D0 U2542 ( .A1(n4101), .A2(n3844), .B1(n3998), .B2(
        \theRegs/completionDataOut[6][40] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[40].enDff/theFlop/N3 ) );
  AO22D0 U2543 ( .A1(n4081), .A2(n3923), .B1(n3998), .B2(
        \theRegs/completionDataOut[6][39] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[39].enDff/theFlop/N3 ) );
  AO22D0 U2544 ( .A1(n3141), .A2(n3896), .B1(n3314), .B2(
        \theRegs/completionDataOut[6][0] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U2545 ( .A1(n4083), .A2(n3996), .B1(n3852), .B2(
        \theRegs/completionDataOut[6][1] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U2546 ( .A1(n4079), .A2(n3945), .B1(n4019), .B2(
        \theRegs/completionDataOut[6][2] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U2547 ( .A1(n4088), .A2(n3945), .B1(n4019), .B2(
        \theRegs/completionDataOut[6][3] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U2548 ( .A1(n4080), .A2(n3896), .B1(n3852), .B2(
        \theRegs/completionDataOut[6][4] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U2549 ( .A1(n4066), .A2(n3945), .B1(n3895), .B2(
        \theRegs/completionDataOut[6][5] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U2550 ( .A1(n3147), .A2(n3896), .B1(n3852), .B2(
        \theRegs/completionDataOut[6][6] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U2551 ( .A1(n4090), .A2(n3945), .B1(n3895), .B2(
        \theRegs/completionDataOut[6][7] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U2552 ( .A1(n4084), .A2(n3945), .B1(n4019), .B2(
        \theRegs/completionDataOut[6][8] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U2553 ( .A1(n4087), .A2(n3945), .B1(n4019), .B2(
        \theRegs/completionDataOut[6][9] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[9].enDff/theFlop/N3 ) );
  AO22D0 U2554 ( .A1(n3151), .A2(n3896), .B1(n3852), .B2(
        \theRegs/completionDataOut[6][10] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[10].enDff/theFlop/N3 ) );
  AO22D0 U2555 ( .A1(n3152), .A2(n3896), .B1(n3852), .B2(
        \theRegs/completionDataOut[6][11] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[11].enDff/theFlop/N3 ) );
  AO22D0 U2556 ( .A1(n3153), .A2(n3473), .B1(n3313), .B2(
        \theRegs/completionDataOut[6][12] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[12].enDff/theFlop/N3 ) );
  AO22D0 U2557 ( .A1(n4055), .A2(n3473), .B1(n3563), .B2(
        \theRegs/completionDataOut[6][13] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[13].enDff/theFlop/N3 ) );
  AO22D0 U2558 ( .A1(n3155), .A2(n3473), .B1(n3313), .B2(
        \theRegs/completionDataOut[6][14] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[14].enDff/theFlop/N3 ) );
  AO22D0 U2559 ( .A1(n4053), .A2(n3473), .B1(n3563), .B2(
        \theRegs/completionDataOut[6][15] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[15].enDff/theFlop/N3 ) );
  AO22D0 U2561 ( .A1(n4049), .A2(n3473), .B1(n3563), .B2(
        \theRegs/completionDataOut[6][16] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[16].enDff/theFlop/N3 ) );
  AO22D0 U2562 ( .A1(n3158), .A2(n3499), .B1(n3600), .B2(
        \theRegs/completionDataOut[6][17] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[17].enDff/theFlop/N3 ) );
  AO22D0 U2564 ( .A1(n4114), .A2(n3709), .B1(n3623), .B2(
        \theRegs/completionDataOut[6][18] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[18].enDff/theFlop/N3 ) );
  AO22D0 U2565 ( .A1(n4044), .A2(n3679), .B1(n3600), .B2(
        \theRegs/completionDataOut[6][19] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[19].enDff/theFlop/N3 ) );
  AO22D0 U2566 ( .A1(n3161), .A2(n3638), .B1(n3438), .B2(
        \theRegs/completionDataOut[6][20] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[20].enDff/theFlop/N3 ) );
  AO22D0 U2567 ( .A1(n3162), .A2(n3638), .B1(n3438), .B2(
        \theRegs/completionDataOut[6][21] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[21].enDff/theFlop/N3 ) );
  AO22D0 U2568 ( .A1(n3163), .A2(n3709), .B1(n3623), .B2(
        \theRegs/completionDataOut[6][22] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[22].enDff/theFlop/N3 ) );
  AO22D0 U2569 ( .A1(n3164), .A2(n3679), .B1(n3600), .B2(
        \theRegs/completionDataOut[6][23] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[23].enDff/theFlop/N3 ) );
  AO22D0 U2572 ( .A1(n3166), .A2(n3679), .B1(n3774), .B2(
        \theRegs/completionDataOut[6][25] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[25].enDff/theFlop/N3 ) );
  AO22D0 U2573 ( .A1(n4102), .A2(n4022), .B1(n3807), .B2(
        \theRegs/completionDataOut[6][49] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[49].enDff/theFlop/N3 ) );
  AO22D0 U2574 ( .A1(n4061), .A2(n3985), .B1(n3807), .B2(
        \theRegs/completionDataOut[6][48] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[48].enDff/theFlop/N3 ) );
  AO22D0 U2575 ( .A1(n3188), .A2(n3679), .B1(n3774), .B2(
        \theRegs/completionDataOut[6][47] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[47].enDff/theFlop/N3 ) );
  AO22D0 U2576 ( .A1(n3170), .A2(n3638), .B1(n3563), .B2(
        \theRegs/completionDataOut[6][29] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[29].enDff/theFlop/N3 ) );
  AO22D0 U2577 ( .A1(n4094), .A2(n3844), .B1(n3998), .B2(
        \theRegs/completionDataOut[6][45] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[45].enDff/theFlop/N3 ) );
  AO22D0 U2578 ( .A1(n4108), .A2(n3749), .B1(n4018), .B2(
        \theRegs/completionDataOut[6][44] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[44].enDff/theFlop/N3 ) );
  AO22D0 U2579 ( .A1(n4100), .A2(n3749), .B1(n4018), .B2(
        \theRegs/completionDataOut[6][43] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[43].enDff/theFlop/N3 ) );
  AO22D0 U2580 ( .A1(n4104), .A2(n3996), .B1(n4019), .B2(
        \theRegs/completionDataOut[6][34] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[34].enDff/theFlop/N3 ) );
  AO22D0 U2581 ( .A1(n3176), .A2(n3896), .B1(n3852), .B2(
        \theRegs/completionDataOut[6][35] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[35].enDff/theFlop/N3 ) );
  AO22D0 U2582 ( .A1(n3177), .A2(n3749), .B1(n4018), .B2(
        \theRegs/completionDataOut[6][36] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[36].enDff/theFlop/N3 ) );
  AO22D0 U2583 ( .A1(n3178), .A2(n3710), .B1(n3970), .B2(
        \theRegs/completionDataOut[6][37] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[37].enDff/theFlop/N3 ) );
  AO22D0 U2584 ( .A1(n3179), .A2(n3749), .B1(n3848), .B2(
        \theRegs/completionDataOut[6][38] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[38].enDff/theFlop/N3 ) );
  AO22D0 U2587 ( .A1(n4098), .A2(n3709), .B1(n3623), .B2(
        \theRegs/completionDataOut[6][24] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[24].enDff/theFlop/N3 ) );
  AO22D0 U2588 ( .A1(n4045), .A2(n3679), .B1(n3600), .B2(
        \theRegs/completionDataOut[6][33] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[33].enDff/theFlop/N3 ) );
  AO22D0 U2589 ( .A1(n3167), .A2(n3915), .B1(n3623), .B2(
        \theRegs/completionDataOut[6][26] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[26].enDff/theFlop/N3 ) );
  AO22D0 U2590 ( .A1(n3168), .A2(n3679), .B1(n3774), .B2(
        \theRegs/completionDataOut[6][27] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[27].enDff/theFlop/N3 ) );
  AO22D0 U2591 ( .A1(n3169), .A2(n3638), .B1(n3563), .B2(
        \theRegs/completionDataOut[6][28] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[28].enDff/theFlop/N3 ) );
  AO22D0 U2592 ( .A1(n3171), .A2(n3499), .B1(n3600), .B2(
        \theRegs/completionDataOut[6][30] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[30].enDff/theFlop/N3 ) );
  AO22D0 U2593 ( .A1(n3172), .A2(n3499), .B1(n3600), .B2(
        \theRegs/completionDataOut[6][31] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[31].enDff/theFlop/N3 ) );
  AO22D0 U2601 ( .A1(n4100), .A2(n3897), .B1(n3388), .B2(
        \theRegs/completionDataOut[2][43] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[43].enDff/theFlop/N3 ) );
  AO22D0 U2602 ( .A1(n4107), .A2(n3994), .B1(n3477), .B2(
        \theRegs/completionDataOut[2][47] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[47].enDff/theFlop/N3 ) );
  AO22D0 U2603 ( .A1(n4076), .A2(n3802), .B1(n3364), .B2(
        \theRegs/completionDataOut[2][46] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[46].enDff/theFlop/N3 ) );
  AO22D0 U2604 ( .A1(n4094), .A2(n3802), .B1(n3364), .B2(
        \theRegs/completionDataOut[2][45] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[45].enDff/theFlop/N3 ) );
  AO22D0 U2605 ( .A1(n4108), .A2(n4025), .B1(n3417), .B2(
        \theRegs/completionDataOut[2][44] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[44].enDff/theFlop/N3 ) );
  AO22D0 U2606 ( .A1(n4072), .A2(n3949), .B1(n3427), .B2(
        \theRegs/completionDataOut[2][36] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[36].enDff/theFlop/N3 ) );
  AO22D0 U2607 ( .A1(n4095), .A2(n3701), .B1(n3361), .B2(
        \theRegs/completionDataOut[2][42] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[42].enDff/theFlop/N3 ) );
  AO22D0 U2608 ( .A1(n4061), .A2(n3949), .B1(n3477), .B2(
        \theRegs/completionDataOut[2][48] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[48].enDff/theFlop/N3 ) );
  AO22D0 U2609 ( .A1(n4101), .A2(n4025), .B1(n3388), .B2(
        \theRegs/completionDataOut[2][40] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[40].enDff/theFlop/N3 ) );
  AO22D0 U2610 ( .A1(n4046), .A2(n3832), .B1(n3761), .B2(
        \theRegs/completionDataOut[2][32] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[32].enDff/theFlop/N3 ) );
  AO22D0 U2611 ( .A1(n4047), .A2(n4001), .B1(n4024), .B2(
        \theRegs/completionDataOut[2][31] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[31].enDff/theFlop/N3 ) );
  AO22D0 U2612 ( .A1(n4051), .A2(n3905), .B1(n3959), .B2(
        \theRegs/completionDataOut[2][30] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[30].enDff/theFlop/N3 ) );
  AO22D0 U2613 ( .A1(n4105), .A2(n3782), .B1(n3686), .B2(
        \theRegs/completionDataOut[2][29] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[29].enDff/theFlop/N3 ) );
  AO22D0 U2614 ( .A1(n4103), .A2(n3782), .B1(n3728), .B2(
        \theRegs/completionDataOut[2][28] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[28].enDff/theFlop/N3 ) );
  AO22D0 U2615 ( .A1(n4109), .A2(n3782), .B1(n3728), .B2(
        \theRegs/completionDataOut[2][27] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[27].enDff/theFlop/N3 ) );
  AO22D0 U2616 ( .A1(n4110), .A2(n3832), .B1(n3761), .B2(
        \theRegs/completionDataOut[2][26] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[26].enDff/theFlop/N3 ) );
  AO22D0 U2617 ( .A1(n3182), .A2(n3339), .B1(n3349), .B2(
        \theRegs/completionDataOut[2][41] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[41].enDff/theFlop/N3 ) );
  AO22D0 U2618 ( .A1(n3165), .A2(n3782), .B1(n3535), .B2(
        \theRegs/completionDataOut[2][24] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[24].enDff/theFlop/N3 ) );
  AO22D0 U2619 ( .A1(n4081), .A2(n3869), .B1(n3351), .B2(
        \theRegs/completionDataOut[2][39] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[39].enDff/theFlop/N3 ) );
  AO22D0 U2620 ( .A1(n3179), .A2(n3701), .B1(n3361), .B2(
        \theRegs/completionDataOut[2][38] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[38].enDff/theFlop/N3 ) );
  AO22D0 U2621 ( .A1(n4077), .A2(n3802), .B1(n3364), .B2(
        \theRegs/completionDataOut[2][37] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[37].enDff/theFlop/N3 ) );
  AO22D0 U2622 ( .A1(n3164), .A2(n3782), .B1(n3535), .B2(
        \theRegs/completionDataOut[2][23] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[23].enDff/theFlop/N3 ) );
  AO22D0 U2623 ( .A1(n4106), .A2(n3802), .B1(n3364), .B2(
        \theRegs/completionDataOut[2][35] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[35].enDff/theFlop/N3 ) );
  AO22D0 U2624 ( .A1(n4104), .A2(n3994), .B1(n3325), .B2(
        \theRegs/completionDataOut[2][34] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[34].enDff/theFlop/N3 ) );
  AO22D0 U2625 ( .A1(n3174), .A2(n3587), .B1(n3325), .B2(
        \theRegs/completionDataOut[2][33] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[33].enDff/theFlop/N3 ) );
  AO22D0 U2626 ( .A1(n3194), .A2(n3785), .B1(n3349), .B2(
        \theRegs/completionDataOut[2][53] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[53].enDff/theFlop/N3 ) );
  AO22D0 U2627 ( .A1(n3193), .A2(n3897), .B1(n3388), .B2(
        \theRegs/completionDataOut[2][52] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[52].enDff/theFlop/N3 ) );
  AO22D0 U2629 ( .A1(n4057), .A2(n3869), .B1(n3381), .B2(
        \theRegs/completionDataOut[2][51] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[51].enDff/theFlop/N3 ) );
  AO22D0 U2630 ( .A1(n4058), .A2(n3949), .B1(n3427), .B2(
        \theRegs/completionDataOut[2][50] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[50].enDff/theFlop/N3 ) );
  AO22D0 U2631 ( .A1(n4102), .A2(n3949), .B1(n3427), .B2(
        \theRegs/completionDataOut[2][49] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[49].enDff/theFlop/N3 ) );
  AO22D0 U2634 ( .A1(n4111), .A2(n3905), .B1(n3959), .B2(
        \theRegs/completionDataOut[2][25] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[25].enDff/theFlop/N3 ) );
  AO22D0 U2635 ( .A1(n3160), .A2(n3340), .B1(n3325), .B2(
        \theRegs/completionDataOut[2][19] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[19].enDff/theFlop/N3 ) );
  AO22D0 U2636 ( .A1(n3141), .A2(n3587), .B1(n3686), .B2(
        \theRegs/completionDataOut[2][0] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U2637 ( .A1(n4083), .A2(n4001), .B1(n4024), .B2(
        \theRegs/completionDataOut[2][1] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U2638 ( .A1(n4079), .A2(n4001), .B1(n4024), .B2(
        \theRegs/completionDataOut[2][2] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U2639 ( .A1(n4088), .A2(n3905), .B1(n3959), .B2(
        \theRegs/completionDataOut[2][3] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U2640 ( .A1(n3145), .A2(n3587), .B1(n3686), .B2(
        \theRegs/completionDataOut[2][4] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U2641 ( .A1(n3146), .A2(n3865), .B1(n3919), .B2(
        \theRegs/completionDataOut[2][5] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U2642 ( .A1(n3147), .A2(n3865), .B1(n3728), .B2(
        \theRegs/completionDataOut[2][6] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U2643 ( .A1(n4090), .A2(n3865), .B1(n3919), .B2(
        \theRegs/completionDataOut[2][7] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U2644 ( .A1(n4084), .A2(n3832), .B1(n3761), .B2(
        \theRegs/completionDataOut[2][8] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U2645 ( .A1(n3150), .A2(n3610), .B1(n3728), .B2(
        \theRegs/completionDataOut[2][9] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[9].enDff/theFlop/N3 ) );
  AO22D0 U2646 ( .A1(n4091), .A2(n3905), .B1(n3959), .B2(
        \theRegs/completionDataOut[2][10] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[10].enDff/theFlop/N3 ) );
  AO22D0 U2647 ( .A1(n3152), .A2(n3587), .B1(n3686), .B2(
        \theRegs/completionDataOut[2][11] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[11].enDff/theFlop/N3 ) );
  AO22D0 U2648 ( .A1(n4056), .A2(n3832), .B1(n3761), .B2(
        \theRegs/completionDataOut[2][12] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[12].enDff/theFlop/N3 ) );
  AO22D0 U2649 ( .A1(n3154), .A2(n3610), .B1(n3728), .B2(
        \theRegs/completionDataOut[2][13] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[13].enDff/theFlop/N3 ) );
  AO22D0 U2650 ( .A1(n4054), .A2(n3865), .B1(n3728), .B2(
        \theRegs/completionDataOut[2][14] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[14].enDff/theFlop/N3 ) );
  AO22D0 U2651 ( .A1(n4053), .A2(n3832), .B1(n3761), .B2(
        \theRegs/completionDataOut[2][15] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[15].enDff/theFlop/N3 ) );
  AO22D0 U2653 ( .A1(n4049), .A2(n4001), .B1(n4024), .B2(
        \theRegs/completionDataOut[2][16] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[16].enDff/theFlop/N3 ) );
  AO22D0 U2654 ( .A1(n4048), .A2(n3905), .B1(n3959), .B2(
        \theRegs/completionDataOut[2][17] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[17].enDff/theFlop/N3 ) );
  AO22D0 U2656 ( .A1(n4114), .A2(n3587), .B1(n3686), .B2(
        \theRegs/completionDataOut[2][18] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[18].enDff/theFlop/N3 ) );
  AO22D0 U2657 ( .A1(n4113), .A2(n3865), .B1(n3919), .B2(
        \theRegs/completionDataOut[2][20] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[20].enDff/theFlop/N3 ) );
  AO22D0 U2658 ( .A1(n4112), .A2(n3832), .B1(n3761), .B2(
        \theRegs/completionDataOut[2][21] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[21].enDff/theFlop/N3 ) );
  AO22D0 U2659 ( .A1(n4092), .A2(n3905), .B1(n3959), .B2(
        \theRegs/completionDataOut[2][22] ), .Z(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[22].enDff/theFlop/N3 ) );
  AO22D0 U2668 ( .A1(n3210), .A2(n3917), .B1(
        \theRegs/completionDataOut[1][69] ), .B2(n3365), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[69].enDff/theFlop/N3 ) );
  AO22D0 U2669 ( .A1(n3210), .A2(n3966), .B1(
        \theRegs/completionDataOut[3][69] ), .B2(n3382), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[69].enDff/theFlop/N3 ) );
  AO22D0 U2670 ( .A1(n3208), .A2(n3966), .B1(n3418), .B2(
        \theRegs/completionDataOut[3][67] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[67].enDff/theFlop/N3 ) );
  AO22D0 U2671 ( .A1(n3209), .A2(n3889), .B1(n3395), .B2(
        \theRegs/completionDataOut[3][68] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[68].enDff/theFlop/N3 ) );
  AO22D0 U2672 ( .A1(n4060), .A2(n3706), .B1(n3365), .B2(
        \theRegs/completionDataOut[1][66] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[66].enDff/theFlop/N3 ) );
  AO22D0 U2673 ( .A1(n3208), .A2(n3706), .B1(n3365), .B2(
        \theRegs/completionDataOut[1][67] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[67].enDff/theFlop/N3 ) );
  AO22D0 U2674 ( .A1(n4059), .A2(n3854), .B1(n3480), .B2(
        \theRegs/completionDataOut[1][68] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[68].enDff/theFlop/N3 ) );
  AO22D0 U2675 ( .A1(n3207), .A2(n3333), .B1(n3318), .B2(
        \theRegs/completionDataOut[3][66] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[66].enDff/theFlop/N3 ) );
  AO22D0 U2676 ( .A1(n4073), .A2(n3898), .B1(n3478), .B2(
        \theRegs/completionDataOut[3][61] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[61].enDff/theFlop/N3 ) );
  AO22D0 U2677 ( .A1(n4064), .A2(n3950), .B1(n3529), .B2(
        \theRegs/completionDataOut[3][65] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[65].enDff/theFlop/N3 ) );
  AO22D0 U2678 ( .A1(n4052), .A2(n3995), .B1(n3590), .B2(
        \theRegs/completionDataOut[3][58] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[58].enDff/theFlop/N3 ) );
  AO22D0 U2679 ( .A1(n3200), .A2(n3833), .B1(n3367), .B2(
        \theRegs/completionDataOut[3][59] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[59].enDff/theFlop/N3 ) );
  AO22D0 U2680 ( .A1(n4078), .A2(n3889), .B1(n3395), .B2(
        \theRegs/completionDataOut[3][60] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[60].enDff/theFlop/N3 ) );
  AO22D0 U2681 ( .A1(n3206), .A2(n3783), .B1(n3357), .B2(
        \theRegs/completionDataOut[1][65] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[65].enDff/theFlop/N3 ) );
  AO22D0 U2682 ( .A1(n3203), .A2(n3748), .B1(n3360), .B2(
        \theRegs/completionDataOut[3][62] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[62].enDff/theFlop/N3 ) );
  AO22D0 U2683 ( .A1(n4071), .A2(n3898), .B1(n3395), .B2(
        \theRegs/completionDataOut[3][63] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[63].enDff/theFlop/N3 ) );
  AO22D0 U2684 ( .A1(n4062), .A2(n3898), .B1(n3478), .B2(
        \theRegs/completionDataOut[3][64] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[64].enDff/theFlop/N3 ) );
  AO22D0 U2685 ( .A1(n4085), .A2(n3898), .B1(n3478), .B2(
        \theRegs/completionDataOut[3][54] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[54].enDff/theFlop/N3 ) );
  AO22D0 U2686 ( .A1(n4074), .A2(n3872), .B1(n3382), .B2(
        \theRegs/completionDataOut[3][55] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[55].enDff/theFlop/N3 ) );
  AO22D0 U2687 ( .A1(n4082), .A2(n3833), .B1(n3367), .B2(
        \theRegs/completionDataOut[3][56] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[56].enDff/theFlop/N3 ) );
  AO22D0 U2688 ( .A1(n4086), .A2(n3995), .B1(n3590), .B2(
        \theRegs/completionDataOut[3][57] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[57].enDff/theFlop/N3 ) );
  AO22D0 U2690 ( .A1(n4074), .A2(n3917), .B1(n3480), .B2(
        \theRegs/completionDataOut[1][55] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[55].enDff/theFlop/N3 ) );
  AO22D0 U2691 ( .A1(n4071), .A2(n3953), .B1(n3510), .B2(
        \theRegs/completionDataOut[1][63] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[63].enDff/theFlop/N3 ) );
  AO22D0 U2692 ( .A1(n4065), .A2(n3990), .B1(n3546), .B2(
        \theRegs/completionDataOut[1][62] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[62].enDff/theFlop/N3 ) );
  AO22D0 U2693 ( .A1(n4073), .A2(n3783), .B1(n3365), .B2(
        \theRegs/completionDataOut[1][61] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[61].enDff/theFlop/N3 ) );
  AO22D0 U2694 ( .A1(n4078), .A2(n3826), .B1(n3389), .B2(
        \theRegs/completionDataOut[1][60] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[60].enDff/theFlop/N3 ) );
  AO22D0 U2695 ( .A1(n4050), .A2(n3953), .B1(n3510), .B2(
        \theRegs/completionDataOut[1][59] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[59].enDff/theFlop/N3 ) );
  AO22D0 U2696 ( .A1(n4052), .A2(n3826), .B1(n3389), .B2(
        \theRegs/completionDataOut[1][58] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[58].enDff/theFlop/N3 ) );
  AO22D0 U2697 ( .A1(n4082), .A2(n3953), .B1(n3510), .B2(
        \theRegs/completionDataOut[1][56] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[56].enDff/theFlop/N3 ) );
  AO22D0 U2698 ( .A1(n4062), .A2(n3917), .B1(n3480), .B2(
        \theRegs/completionDataOut[1][64] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[64].enDff/theFlop/N3 ) );
  AO22D0 U2699 ( .A1(n4085), .A2(n3990), .B1(n3546), .B2(
        \theRegs/completionDataOut[1][54] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[54].enDff/theFlop/N3 ) );
  AO22D0 U2700 ( .A1(n3198), .A2(n3336), .B1(n3357), .B2(
        \theRegs/completionDataOut[1][57] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[57].enDff/theFlop/N3 ) );
  AO22D0 U2702 ( .A1(n3205), .A2(n3391), .B1(n3729), .B2(
        \theRegs/completionDataOut[5][64] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[64].enDff/theFlop/N3 ) );
  AO22D0 U2703 ( .A1(n4059), .A2(n3700), .B1(n3944), .B2(
        \theRegs/completionDataOut[5][68] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[68].enDff/theFlop/N3 ) );
  AO22D0 U2704 ( .A1(n3206), .A2(n3483), .B1(n3868), .B2(
        \theRegs/completionDataOut[5][65] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[65].enDff/theFlop/N3 ) );
  AO22D0 U2705 ( .A1(n3207), .A2(n3380), .B1(n3687), .B2(
        \theRegs/completionDataOut[5][66] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[66].enDff/theFlop/N3 ) );
  AO22D0 U2706 ( .A1(n3196), .A2(n3380), .B1(n3687), .B2(
        \theRegs/completionDataOut[5][55] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[55].enDff/theFlop/N3 ) );
  AO22D0 U2707 ( .A1(n3195), .A2(n3391), .B1(n3729), .B2(
        \theRegs/completionDataOut[5][54] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[54].enDff/theFlop/N3 ) );
  AO22D0 U2708 ( .A1(n4078), .A2(n3627), .B1(n3964), .B2(
        \theRegs/completionDataOut[5][60] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[60].enDff/theFlop/N3 ) );
  AO22D0 U2709 ( .A1(n3202), .A2(n3380), .B1(n3687), .B2(
        \theRegs/completionDataOut[5][61] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[61].enDff/theFlop/N3 ) );
  AO22D0 U2710 ( .A1(n4065), .A2(n3700), .B1(n3944), .B2(
        \theRegs/completionDataOut[5][62] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[62].enDff/theFlop/N3 ) );
  AO22D0 U2711 ( .A1(n3208), .A2(n3423), .B1(n3729), .B2(
        \theRegs/completionDataOut[5][67] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[67].enDff/theFlop/N3 ) );
  AO22D0 U2712 ( .A1(n4068), .A2(n3700), .B1(
        \theRegs/completionDataOut[5][69] ), .B2(n3964), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[69].enDff/theFlop/N3 ) );
  AO22D0 U2713 ( .A1(n4086), .A2(n3433), .B1(n3742), .B2(
        \theRegs/completionDataOut[5][57] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[57].enDff/theFlop/N3 ) );
  AO22D0 U2714 ( .A1(n3197), .A2(n3380), .B1(n3338), .B2(
        \theRegs/completionDataOut[5][56] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[56].enDff/theFlop/N3 ) );
  AO22D0 U2715 ( .A1(n4050), .A2(n3433), .B1(n3742), .B2(
        \theRegs/completionDataOut[5][59] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[59].enDff/theFlop/N3 ) );
  AO22D0 U2716 ( .A1(n3199), .A2(n3391), .B1(n3729), .B2(
        \theRegs/completionDataOut[5][58] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[58].enDff/theFlop/N3 ) );
  AO22D0 U2717 ( .A1(n4071), .A2(n3700), .B1(n3944), .B2(
        \theRegs/completionDataOut[5][63] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[63].enDff/theFlop/N3 ) );
  AO22D0 U2719 ( .A1(n4102), .A2(n3784), .B1(n3944), .B2(
        \theRegs/completionDataOut[5][49] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[49].enDff/theFlop/N3 ) );
  AO22D0 U2720 ( .A1(n3146), .A2(n4002), .B1(n4023), .B2(
        \theRegs/completionDataOut[3][5] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U2721 ( .A1(n4070), .A2(n3483), .B1(n3868), .B2(
        \theRegs/completionDataOut[5][53] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[53].enDff/theFlop/N3 ) );
  AO22D0 U2722 ( .A1(n4057), .A2(n3423), .B1(n3729), .B2(
        \theRegs/completionDataOut[5][51] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[51].enDff/theFlop/N3 ) );
  AO22D0 U2723 ( .A1(n4107), .A2(n3872), .B1(n3360), .B2(
        \theRegs/completionDataOut[3][47] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[47].enDff/theFlop/N3 ) );
  AO22D0 U2724 ( .A1(n4061), .A2(n4026), .B1(n3395), .B2(
        \theRegs/completionDataOut[3][48] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[48].enDff/theFlop/N3 ) );
  AO22D0 U2725 ( .A1(n4102), .A2(n3898), .B1(n3478), .B2(
        \theRegs/completionDataOut[3][49] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[49].enDff/theFlop/N3 ) );
  AO22D0 U2726 ( .A1(n3191), .A2(n3872), .B1(n3360), .B2(
        \theRegs/completionDataOut[3][50] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[50].enDff/theFlop/N3 ) );
  AO22D0 U2727 ( .A1(n4057), .A2(n3872), .B1(n3382), .B2(
        \theRegs/completionDataOut[3][51] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[51].enDff/theFlop/N3 ) );
  AO22D0 U2728 ( .A1(n4067), .A2(n3950), .B1(n3529), .B2(
        \theRegs/completionDataOut[3][52] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[52].enDff/theFlop/N3 ) );
  AO22D0 U2729 ( .A1(n4070), .A2(n3833), .B1(n3418), .B2(
        \theRegs/completionDataOut[3][53] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[53].enDff/theFlop/N3 ) );
  AO22D0 U2731 ( .A1(n3193), .A2(n3433), .B1(n3742), .B2(
        \theRegs/completionDataOut[5][52] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[52].enDff/theFlop/N3 ) );
  AO22D0 U2733 ( .A1(n4102), .A2(n3953), .B1(n3510), .B2(
        \theRegs/completionDataOut[1][49] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[49].enDff/theFlop/N3 ) );
  AO22D0 U2734 ( .A1(n4058), .A2(n3854), .B1(n3480), .B2(
        \theRegs/completionDataOut[1][50] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[50].enDff/theFlop/N3 ) );
  AO22D0 U2735 ( .A1(n3192), .A2(n3783), .B1(n3384), .B2(
        \theRegs/completionDataOut[1][51] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[51].enDff/theFlop/N3 ) );
  AO22D0 U2736 ( .A1(n3193), .A2(n3990), .B1(n3546), .B2(
        \theRegs/completionDataOut[1][52] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[52].enDff/theFlop/N3 ) );
  AO22D0 U2737 ( .A1(n4070), .A2(n3706), .B1(n3420), .B2(
        \theRegs/completionDataOut[1][53] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[53].enDff/theFlop/N3 ) );
  AO22D0 U2739 ( .A1(n4058), .A2(n3784), .B1(n3997), .B2(
        \theRegs/completionDataOut[5][50] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[50].enDff/theFlop/N3 ) );
  AO22D0 U2740 ( .A1(n4107), .A2(n3433), .B1(n3742), .B2(
        \theRegs/completionDataOut[5][47] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[47].enDff/theFlop/N3 ) );
  AO22D0 U2741 ( .A1(n3189), .A2(n3380), .B1(n3687), .B2(
        \theRegs/completionDataOut[5][48] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[48].enDff/theFlop/N3 ) );
  AO22D0 U2742 ( .A1(n4101), .A2(n3950), .B1(n3529), .B2(
        \theRegs/completionDataOut[3][40] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[40].enDff/theFlop/N3 ) );
  AO22D0 U2743 ( .A1(n4061), .A2(n3953), .B1(n3510), .B2(
        \theRegs/completionDataOut[1][48] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[48].enDff/theFlop/N3 ) );
  AO22D0 U2744 ( .A1(n4097), .A2(n3872), .B1(n3382), .B2(
        \theRegs/completionDataOut[3][41] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[41].enDff/theFlop/N3 ) );
  AO22D0 U2745 ( .A1(n4095), .A2(n3966), .B1(n3395), .B2(
        \theRegs/completionDataOut[3][42] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[42].enDff/theFlop/N3 ) );
  AO22D0 U2746 ( .A1(n3184), .A2(n3333), .B1(n3360), .B2(
        \theRegs/completionDataOut[3][43] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[43].enDff/theFlop/N3 ) );
  AO22D0 U2747 ( .A1(n4108), .A2(n3966), .B1(n3418), .B2(
        \theRegs/completionDataOut[3][44] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[44].enDff/theFlop/N3 ) );
  AO22D0 U2748 ( .A1(n4094), .A2(n3966), .B1(n3395), .B2(
        \theRegs/completionDataOut[3][45] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[45].enDff/theFlop/N3 ) );
  AO22D0 U2749 ( .A1(n3187), .A2(n3833), .B1(n3367), .B2(
        \theRegs/completionDataOut[3][46] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[46].enDff/theFlop/N3 ) );
  AO22D0 U2750 ( .A1(n4098), .A2(n3575), .B1(n3702), .B2(
        \theRegs/completionDataOut[5][24] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[24].enDff/theFlop/N3 ) );
  AO22D0 U2751 ( .A1(n3141), .A2(n3322), .B1(n3337), .B2(
        \theRegs/completionDataOut[5][0] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U2752 ( .A1(n3143), .A2(n3870), .B1(n3924), .B2(
        \theRegs/completionDataOut[5][2] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U2753 ( .A1(n4088), .A2(n3904), .B1(n3957), .B2(
        \theRegs/completionDataOut[5][3] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U2754 ( .A1(n4080), .A2(n3870), .B1(n3924), .B2(
        \theRegs/completionDataOut[5][4] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U2755 ( .A1(n4066), .A2(n3999), .B1(n4021), .B2(
        \theRegs/completionDataOut[5][5] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U2756 ( .A1(n4089), .A2(n3759), .B1(n3805), .B2(
        \theRegs/completionDataOut[5][6] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U2757 ( .A1(n4090), .A2(n3904), .B1(n3957), .B2(
        \theRegs/completionDataOut[5][7] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U2758 ( .A1(n3149), .A2(n3575), .B1(n3702), .B2(
        \theRegs/completionDataOut[5][8] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U2759 ( .A1(n3150), .A2(n3322), .B1(n3337), .B2(
        \theRegs/completionDataOut[5][9] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[9].enDff/theFlop/N3 ) );
  AO22D0 U2760 ( .A1(n4091), .A2(n3322), .B1(n3337), .B2(
        \theRegs/completionDataOut[5][10] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[10].enDff/theFlop/N3 ) );
  AO22D0 U2761 ( .A1(n4099), .A2(n3999), .B1(n4021), .B2(
        \theRegs/completionDataOut[5][11] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[11].enDff/theFlop/N3 ) );
  AO22D0 U2762 ( .A1(n4056), .A2(n3759), .B1(n3805), .B2(
        \theRegs/completionDataOut[5][12] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[12].enDff/theFlop/N3 ) );
  AO22D0 U2763 ( .A1(n4055), .A2(n3999), .B1(n4021), .B2(
        \theRegs/completionDataOut[5][13] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[13].enDff/theFlop/N3 ) );
  AO22D0 U2764 ( .A1(n4054), .A2(n3759), .B1(n3805), .B2(
        \theRegs/completionDataOut[5][14] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[14].enDff/theFlop/N3 ) );
  AO22D0 U2765 ( .A1(n4053), .A2(n3575), .B1(n3702), .B2(
        \theRegs/completionDataOut[5][15] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[15].enDff/theFlop/N3 ) );
  AO22D0 U2766 ( .A1(n4049), .A2(n3575), .B1(n3702), .B2(
        \theRegs/completionDataOut[5][16] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[16].enDff/theFlop/N3 ) );
  AO22D0 U2767 ( .A1(n4048), .A2(n3904), .B1(n3957), .B2(
        \theRegs/completionDataOut[5][17] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[17].enDff/theFlop/N3 ) );
  AO22D0 U2768 ( .A1(n4114), .A2(n3575), .B1(n3702), .B2(
        \theRegs/completionDataOut[5][18] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[18].enDff/theFlop/N3 ) );
  AO22D0 U2769 ( .A1(n4044), .A2(n3904), .B1(n3957), .B2(
        \theRegs/completionDataOut[5][19] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[19].enDff/theFlop/N3 ) );
  AO22D0 U2770 ( .A1(n4113), .A2(n3759), .B1(n3805), .B2(
        \theRegs/completionDataOut[5][20] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[20].enDff/theFlop/N3 ) );
  AO22D0 U2771 ( .A1(n4112), .A2(n3575), .B1(n3702), .B2(
        \theRegs/completionDataOut[5][21] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[21].enDff/theFlop/N3 ) );
  AO22D0 U2772 ( .A1(n3163), .A2(n3640), .B1(n3786), .B2(
        \theRegs/completionDataOut[5][22] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[22].enDff/theFlop/N3 ) );
  AO22D0 U2773 ( .A1(n4093), .A2(n3870), .B1(n3924), .B2(
        \theRegs/completionDataOut[5][23] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[23].enDff/theFlop/N3 ) );
  AO22D0 U2774 ( .A1(n4111), .A2(n3904), .B1(n3957), .B2(
        \theRegs/completionDataOut[5][25] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[25].enDff/theFlop/N3 ) );
  AO22D0 U2775 ( .A1(n4110), .A2(n3640), .B1(n3786), .B2(
        \theRegs/completionDataOut[5][26] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[26].enDff/theFlop/N3 ) );
  AO22D0 U2776 ( .A1(n4109), .A2(n3759), .B1(n3805), .B2(
        \theRegs/completionDataOut[5][27] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[27].enDff/theFlop/N3 ) );
  AO22D0 U2777 ( .A1(n4103), .A2(n3904), .B1(n3957), .B2(
        \theRegs/completionDataOut[5][28] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[28].enDff/theFlop/N3 ) );
  AO22D0 U2778 ( .A1(n4105), .A2(n3999), .B1(n4021), .B2(
        \theRegs/completionDataOut[5][29] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[29].enDff/theFlop/N3 ) );
  AO22D0 U2779 ( .A1(n4051), .A2(n3811), .B1(n3997), .B2(
        \theRegs/completionDataOut[5][30] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[30].enDff/theFlop/N3 ) );
  AO22D0 U2780 ( .A1(n4047), .A2(n3627), .B1(n3964), .B2(
        \theRegs/completionDataOut[5][31] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[31].enDff/theFlop/N3 ) );
  AO22D0 U2781 ( .A1(n4046), .A2(n3627), .B1(n3888), .B2(
        \theRegs/completionDataOut[5][32] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[32].enDff/theFlop/N3 ) );
  AO22D0 U2782 ( .A1(n4045), .A2(n3391), .B1(n3729), .B2(
        \theRegs/completionDataOut[5][33] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[33].enDff/theFlop/N3 ) );
  AO22D0 U2784 ( .A1(n4104), .A2(n3811), .B1(n4016), .B2(
        \theRegs/completionDataOut[5][34] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[34].enDff/theFlop/N3 ) );
  AO22D0 U2785 ( .A1(n4106), .A2(n3567), .B1(n3888), .B2(
        \theRegs/completionDataOut[5][35] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[35].enDff/theFlop/N3 ) );
  AO22D0 U2787 ( .A1(n3177), .A2(n3627), .B1(n3964), .B2(
        \theRegs/completionDataOut[5][36] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[36].enDff/theFlop/N3 ) );
  AO22D0 U2788 ( .A1(n4077), .A2(n3483), .B1(n3868), .B2(
        \theRegs/completionDataOut[5][37] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[37].enDff/theFlop/N3 ) );
  AO22D0 U2789 ( .A1(n3179), .A2(n3380), .B1(n3687), .B2(
        \theRegs/completionDataOut[5][38] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[38].enDff/theFlop/N3 ) );
  AO22D0 U2790 ( .A1(n4081), .A2(n3811), .B1(n3894), .B2(
        \theRegs/completionDataOut[5][39] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[39].enDff/theFlop/N3 ) );
  AO22D0 U2791 ( .A1(n4101), .A2(n3784), .B1(n3894), .B2(
        \theRegs/completionDataOut[5][40] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[40].enDff/theFlop/N3 ) );
  AO22D0 U2792 ( .A1(n4097), .A2(n3567), .B1(n4016), .B2(
        \theRegs/completionDataOut[5][41] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[41].enDff/theFlop/N3 ) );
  AO22D0 U2793 ( .A1(n4095), .A2(n3700), .B1(n3944), .B2(
        \theRegs/completionDataOut[5][42] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[42].enDff/theFlop/N3 ) );
  AO22D0 U2794 ( .A1(n4100), .A2(n3627), .B1(n3964), .B2(
        \theRegs/completionDataOut[5][43] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[43].enDff/theFlop/N3 ) );
  AO22D0 U2795 ( .A1(n4108), .A2(n3423), .B1(n3687), .B2(
        \theRegs/completionDataOut[5][44] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[44].enDff/theFlop/N3 ) );
  AO22D0 U2796 ( .A1(n4094), .A2(n3811), .B1(n4016), .B2(
        \theRegs/completionDataOut[5][45] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[45].enDff/theFlop/N3 ) );
  AO22D0 U2797 ( .A1(n4076), .A2(n3811), .B1(n4016), .B2(
        \theRegs/completionDataOut[5][46] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[46].enDff/theFlop/N3 ) );
  AO22D0 U2801 ( .A1(n3142), .A2(n3759), .B1(n3805), .B2(
        \theRegs/completionDataOut[5][1] ), .Z(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U2809 ( .A1(n4107), .A2(n3706), .B1(n3365), .B2(
        \theRegs/completionDataOut[1][47] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[47].enDff/theFlop/N3 ) );
  AO22D0 U2810 ( .A1(n3187), .A2(n3783), .B1(n3384), .B2(
        \theRegs/completionDataOut[1][46] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[46].enDff/theFlop/N3 ) );
  AO22D0 U2811 ( .A1(n4094), .A2(n3826), .B1(n3389), .B2(
        \theRegs/completionDataOut[1][45] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[45].enDff/theFlop/N3 ) );
  AO22D0 U2812 ( .A1(n4108), .A2(n3826), .B1(n3389), .B2(
        \theRegs/completionDataOut[1][44] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[44].enDff/theFlop/N3 ) );
  AO22D0 U2813 ( .A1(n4100), .A2(n3953), .B1(n3510), .B2(
        \theRegs/completionDataOut[1][43] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[43].enDff/theFlop/N3 ) );
  AO22D0 U2814 ( .A1(n4095), .A2(n3990), .B1(n3546), .B2(
        \theRegs/completionDataOut[1][42] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[42].enDff/theFlop/N3 ) );
  AO22D0 U2815 ( .A1(n4097), .A2(n3336), .B1(n3357), .B2(
        \theRegs/completionDataOut[1][41] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[41].enDff/theFlop/N3 ) );
  AO22D0 U2816 ( .A1(n4101), .A2(n3854), .B1(n3430), .B2(
        \theRegs/completionDataOut[1][40] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[40].enDff/theFlop/N3 ) );
  AO22D0 U2817 ( .A1(n4081), .A2(n3826), .B1(n3389), .B2(
        \theRegs/completionDataOut[1][39] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[39].enDff/theFlop/N3 ) );
  AO22D0 U2818 ( .A1(n4063), .A2(n3826), .B1(n3389), .B2(
        \theRegs/completionDataOut[1][38] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[38].enDff/theFlop/N3 ) );
  AO22D0 U2819 ( .A1(n4077), .A2(n3706), .B1(n3365), .B2(
        \theRegs/completionDataOut[1][37] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[37].enDff/theFlop/N3 ) );
  AO22D0 U2820 ( .A1(n3177), .A2(n3917), .B1(n3480), .B2(
        \theRegs/completionDataOut[1][36] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[36].enDff/theFlop/N3 ) );
  AO22D0 U2822 ( .A1(n4106), .A2(n3854), .B1(n3430), .B2(
        \theRegs/completionDataOut[1][35] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[35].enDff/theFlop/N3 ) );
  AO22D0 U2823 ( .A1(n4104), .A2(n3917), .B1(n3484), .B2(
        \theRegs/completionDataOut[1][34] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[34].enDff/theFlop/N3 ) );
  AO22D0 U2825 ( .A1(n4045), .A2(n3954), .B1(n3665), .B2(
        \theRegs/completionDataOut[1][33] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[33].enDff/theFlop/N3 ) );
  AO22D0 U2826 ( .A1(n4046), .A2(n3954), .B1(n3606), .B2(
        \theRegs/completionDataOut[1][32] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[32].enDff/theFlop/N3 ) );
  AO22D0 U2827 ( .A1(n4047), .A2(n3875), .B1(n3506), .B2(
        \theRegs/completionDataOut[1][31] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[31].enDff/theFlop/N3 ) );
  AO22D0 U2828 ( .A1(n4051), .A2(n3918), .B1(n3484), .B2(
        \theRegs/completionDataOut[1][30] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[30].enDff/theFlop/N3 ) );
  AO22D0 U2829 ( .A1(n4105), .A2(n3763), .B1(n3413), .B2(
        \theRegs/completionDataOut[1][29] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[29].enDff/theFlop/N3 ) );
  AO22D0 U2830 ( .A1(n4103), .A2(n3828), .B1(n3453), .B2(
        \theRegs/completionDataOut[1][28] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[28].enDff/theFlop/N3 ) );
  AO22D0 U2831 ( .A1(n4109), .A2(n3918), .B1(n3484), .B2(
        \theRegs/completionDataOut[1][27] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[27].enDff/theFlop/N3 ) );
  AO22D0 U2832 ( .A1(n4110), .A2(n3828), .B1(n3393), .B2(
        \theRegs/completionDataOut[1][26] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[26].enDff/theFlop/N3 ) );
  AO22D0 U2833 ( .A1(n4111), .A2(n3335), .B1(n3393), .B2(
        \theRegs/completionDataOut[1][25] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[25].enDff/theFlop/N3 ) );
  AO22D0 U2834 ( .A1(n4098), .A2(n3918), .B1(n3484), .B2(
        \theRegs/completionDataOut[1][24] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[24].enDff/theFlop/N3 ) );
  AO22D0 U2835 ( .A1(n4093), .A2(n3875), .B1(n3506), .B2(
        \theRegs/completionDataOut[1][23] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[23].enDff/theFlop/N3 ) );
  AO22D0 U2836 ( .A1(n4092), .A2(n3954), .B1(n3665), .B2(
        \theRegs/completionDataOut[1][22] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[22].enDff/theFlop/N3 ) );
  AO22D0 U2837 ( .A1(n4112), .A2(n3828), .B1(n3453), .B2(
        \theRegs/completionDataOut[1][21] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[21].enDff/theFlop/N3 ) );
  AO22D0 U2838 ( .A1(n4113), .A2(n3763), .B1(n3453), .B2(
        \theRegs/completionDataOut[1][20] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[20].enDff/theFlop/N3 ) );
  AO22D0 U2839 ( .A1(n4044), .A2(n3991), .B1(n3665), .B2(
        \theRegs/completionDataOut[1][19] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[19].enDff/theFlop/N3 ) );
  AO22D0 U2840 ( .A1(n4114), .A2(n3875), .B1(n3548), .B2(
        \theRegs/completionDataOut[1][18] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[18].enDff/theFlop/N3 ) );
  AO22D0 U2842 ( .A1(n4048), .A2(n3991), .B1(n3506), .B2(
        \theRegs/completionDataOut[1][17] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[17].enDff/theFlop/N3 ) );
  AO22D0 U2843 ( .A1(n4049), .A2(n3763), .B1(n3413), .B2(
        \theRegs/completionDataOut[1][16] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[16].enDff/theFlop/N3 ) );
  AO22D0 U2846 ( .A1(n4053), .A2(n3918), .B1(n3484), .B2(
        \theRegs/completionDataOut[1][15] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[15].enDff/theFlop/N3 ) );
  AO22D0 U2847 ( .A1(n4054), .A2(n3828), .B1(n3413), .B2(
        \theRegs/completionDataOut[1][14] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[14].enDff/theFlop/N3 ) );
  AO22D0 U2848 ( .A1(n4055), .A2(n3335), .B1(n3393), .B2(
        \theRegs/completionDataOut[1][13] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[13].enDff/theFlop/N3 ) );
  AO22D0 U2849 ( .A1(n4056), .A2(n3875), .B1(n3506), .B2(
        \theRegs/completionDataOut[1][12] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[12].enDff/theFlop/N3 ) );
  AO22D0 U2850 ( .A1(n4099), .A2(n3875), .B1(n3548), .B2(
        \theRegs/completionDataOut[1][11] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[11].enDff/theFlop/N3 ) );
  AO22D0 U2851 ( .A1(n4091), .A2(n3335), .B1(n3393), .B2(
        \theRegs/completionDataOut[1][10] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[10].enDff/theFlop/N3 ) );
  AO22D0 U2852 ( .A1(n4087), .A2(n3954), .B1(n3606), .B2(
        \theRegs/completionDataOut[1][9] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[9].enDff/theFlop/N3 ) );
  AO22D0 U2853 ( .A1(n3149), .A2(n3763), .B1(n3413), .B2(
        \theRegs/completionDataOut[1][8] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U2854 ( .A1(n4090), .A2(n3954), .B1(n3665), .B2(
        \theRegs/completionDataOut[1][7] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U2855 ( .A1(n4089), .A2(n3918), .B1(n3484), .B2(
        \theRegs/completionDataOut[1][6] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U2856 ( .A1(n4066), .A2(n3991), .B1(n3506), .B2(
        \theRegs/completionDataOut[1][5] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U2857 ( .A1(n4080), .A2(n3991), .B1(n3506), .B2(
        \theRegs/completionDataOut[1][4] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U2858 ( .A1(n3144), .A2(n3875), .B1(n3548), .B2(
        \theRegs/completionDataOut[1][3] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U2859 ( .A1(n4079), .A2(n3954), .B1(n3665), .B2(
        \theRegs/completionDataOut[1][2] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U2860 ( .A1(n3142), .A2(n3763), .B1(n3413), .B2(
        \theRegs/completionDataOut[1][1] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U2861 ( .A1(n4075), .A2(n3763), .B1(n3413), .B2(
        \theRegs/completionDataOut[1][0] ), .Z(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U2869 ( .A1(n3141), .A2(n3334), .B1(n3574), .B2(
        \theRegs/completionDataOut[3][0] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U2870 ( .A1(n4083), .A2(n4002), .B1(n4023), .B2(
        \theRegs/completionDataOut[3][1] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U2871 ( .A1(n3143), .A2(n3730), .B1(n3574), .B2(
        \theRegs/completionDataOut[3][2] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U2872 ( .A1(n3144), .A2(n3662), .B1(n3624), .B2(
        \theRegs/completionDataOut[3][3] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U2873 ( .A1(n3145), .A2(n3730), .B1(n3319), .B2(
        \theRegs/completionDataOut[3][4] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U2874 ( .A1(n4081), .A2(n3748), .B1(n3360), .B2(
        \theRegs/completionDataOut[3][39] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[39].enDff/theFlop/N3 ) );
  AO22D0 U2875 ( .A1(n4063), .A2(n3833), .B1(n3367), .B2(
        \theRegs/completionDataOut[3][38] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[38].enDff/theFlop/N3 ) );
  AO22D0 U2876 ( .A1(n4077), .A2(n3898), .B1(n3478), .B2(
        \theRegs/completionDataOut[3][37] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[37].enDff/theFlop/N3 ) );
  AO22D0 U2877 ( .A1(n4072), .A2(n3995), .B1(n3590), .B2(
        \theRegs/completionDataOut[3][36] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[36].enDff/theFlop/N3 ) );
  AO22D0 U2879 ( .A1(n4106), .A2(n3833), .B1(n3367), .B2(
        \theRegs/completionDataOut[3][35] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[35].enDff/theFlop/N3 ) );
  AO22D0 U2880 ( .A1(n4104), .A2(n3995), .B1(n3428), .B2(
        \theRegs/completionDataOut[3][34] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[34].enDff/theFlop/N3 ) );
  AO22D0 U2882 ( .A1(n4045), .A2(n3995), .B1(n3428), .B2(
        \theRegs/completionDataOut[3][33] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[33].enDff/theFlop/N3 ) );
  AO22D0 U2883 ( .A1(n4046), .A2(n3950), .B1(n3529), .B2(
        \theRegs/completionDataOut[3][32] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[32].enDff/theFlop/N3 ) );
  AO22D0 U2884 ( .A1(n4047), .A2(n3334), .B1(n3574), .B2(
        \theRegs/completionDataOut[3][31] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[31].enDff/theFlop/N3 ) );
  AO22D0 U2885 ( .A1(n4051), .A2(n3906), .B1(n3958), .B2(
        \theRegs/completionDataOut[3][30] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[30].enDff/theFlop/N3 ) );
  AO22D0 U2886 ( .A1(n4105), .A2(n4002), .B1(n4023), .B2(
        \theRegs/completionDataOut[3][29] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[29].enDff/theFlop/N3 ) );
  AO22D0 U2887 ( .A1(n4103), .A2(n3906), .B1(n3958), .B2(
        \theRegs/completionDataOut[3][28] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[28].enDff/theFlop/N3 ) );
  AO22D0 U2888 ( .A1(n4109), .A2(n3867), .B1(n3922), .B2(
        \theRegs/completionDataOut[3][27] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[27].enDff/theFlop/N3 ) );
  AO22D0 U2889 ( .A1(n4110), .A2(n4002), .B1(n4023), .B2(
        \theRegs/completionDataOut[3][26] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[26].enDff/theFlop/N3 ) );
  AO22D0 U2890 ( .A1(n4111), .A2(n3906), .B1(n3958), .B2(
        \theRegs/completionDataOut[3][25] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[25].enDff/theFlop/N3 ) );
  AO22D0 U2891 ( .A1(n4098), .A2(n3758), .B1(n3804), .B2(
        \theRegs/completionDataOut[3][24] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[24].enDff/theFlop/N3 ) );
  AO22D0 U2892 ( .A1(n4093), .A2(n3758), .B1(n3804), .B2(
        \theRegs/completionDataOut[3][23] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[23].enDff/theFlop/N3 ) );
  AO22D0 U2893 ( .A1(n3163), .A2(n3662), .B1(n3624), .B2(
        \theRegs/completionDataOut[3][22] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[22].enDff/theFlop/N3 ) );
  AO22D0 U2894 ( .A1(n4112), .A2(n3758), .B1(n3804), .B2(
        \theRegs/completionDataOut[3][21] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[21].enDff/theFlop/N3 ) );
  AO22D0 U2895 ( .A1(n4113), .A2(n3662), .B1(n3624), .B2(
        \theRegs/completionDataOut[3][20] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[20].enDff/theFlop/N3 ) );
  AO22D0 U2896 ( .A1(n4044), .A2(n3906), .B1(n3958), .B2(
        \theRegs/completionDataOut[3][19] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[19].enDff/theFlop/N3 ) );
  AO22D0 U2897 ( .A1(n4114), .A2(n3730), .B1(n3319), .B2(
        \theRegs/completionDataOut[3][18] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[18].enDff/theFlop/N3 ) );
  AO22D0 U2899 ( .A1(n4048), .A2(n3758), .B1(n3804), .B2(
        \theRegs/completionDataOut[3][17] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[17].enDff/theFlop/N3 ) );
  AO22D0 U2900 ( .A1(n4049), .A2(n3730), .B1(n3319), .B2(
        \theRegs/completionDataOut[3][16] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[16].enDff/theFlop/N3 ) );
  AO22D0 U2903 ( .A1(n4053), .A2(n3662), .B1(n3624), .B2(
        \theRegs/completionDataOut[3][15] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[15].enDff/theFlop/N3 ) );
  AO22D0 U2904 ( .A1(n4054), .A2(n3867), .B1(n3922), .B2(
        \theRegs/completionDataOut[3][14] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[14].enDff/theFlop/N3 ) );
  AO22D0 U2905 ( .A1(n4055), .A2(n3906), .B1(n3958), .B2(
        \theRegs/completionDataOut[3][13] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[13].enDff/theFlop/N3 ) );
  AO22D0 U2906 ( .A1(n4056), .A2(n3334), .B1(n3574), .B2(
        \theRegs/completionDataOut[3][12] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[12].enDff/theFlop/N3 ) );
  AO22D0 U2907 ( .A1(n4099), .A2(n3758), .B1(n3804), .B2(
        \theRegs/completionDataOut[3][11] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[11].enDff/theFlop/N3 ) );
  AO22D0 U2908 ( .A1(n4091), .A2(n3662), .B1(n3624), .B2(
        \theRegs/completionDataOut[3][10] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[10].enDff/theFlop/N3 ) );
  AO22D0 U2909 ( .A1(n4087), .A2(n3867), .B1(n3922), .B2(
        \theRegs/completionDataOut[3][9] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[9].enDff/theFlop/N3 ) );
  AO22D0 U2910 ( .A1(n4084), .A2(n3758), .B1(n3804), .B2(
        \theRegs/completionDataOut[3][8] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U2911 ( .A1(n4090), .A2(n3906), .B1(n3958), .B2(
        \theRegs/completionDataOut[3][7] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U2912 ( .A1(n4089), .A2(n3662), .B1(n3624), .B2(
        \theRegs/completionDataOut[3][6] ), .Z(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U2920 ( .A1(n4068), .A2(n3376), .B1(
        \theRegs/completionDataOut[7][69] ), .B2(n3652), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[69].enDff/theFlop/N3 ) );
  AO22D0 U2921 ( .A1(n3555), .A2(n3208), .B1(n3635), .B2(
        \theRegs/completionDataOut[7][67] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[67].enDff/theFlop/N3 ) );
  AO22D0 U2922 ( .A1(n3740), .A2(n3209), .B1(n3797), .B2(
        \theRegs/completionDataOut[7][68] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[68].enDff/theFlop/N3 ) );
  AO22D0 U2923 ( .A1(n3722), .A2(n3207), .B1(n3775), .B2(
        \theRegs/completionDataOut[7][66] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[66].enDff/theFlop/N3 ) );
  AO22D0 U2924 ( .A1(n3602), .A2(n3197), .B1(n3735), .B2(
        \theRegs/completionDataOut[7][56] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[56].enDff/theFlop/N3 ) );
  AO22D0 U2925 ( .A1(n3331), .A2(n3195), .B1(n3316), .B2(
        \theRegs/completionDataOut[7][54] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[54].enDff/theFlop/N3 ) );
  AO22D0 U2926 ( .A1(n3536), .A2(n3196), .B1(n3735), .B2(
        \theRegs/completionDataOut[7][55] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[55].enDff/theFlop/N3 ) );
  AO22D0 U2927 ( .A1(n3376), .A2(n3206), .B1(n3491), .B2(
        \theRegs/completionDataOut[7][65] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[65].enDff/theFlop/N3 ) );
  AO22D0 U2928 ( .A1(n3740), .A2(n4062), .B1(n3911), .B2(
        \theRegs/completionDataOut[7][64] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[64].enDff/theFlop/N3 ) );
  AO22D0 U2929 ( .A1(n3332), .A2(n3204), .B1(n3317), .B2(
        \theRegs/completionDataOut[7][63] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[63].enDff/theFlop/N3 ) );
  AO22D0 U2930 ( .A1(n3332), .A2(n3203), .B1(n3317), .B2(
        \theRegs/completionDataOut[7][62] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[62].enDff/theFlop/N3 ) );
  AO22D0 U2931 ( .A1(n3376), .A2(n3202), .B1(n3491), .B2(
        \theRegs/completionDataOut[7][61] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[61].enDff/theFlop/N3 ) );
  AO22D0 U2932 ( .A1(n3376), .A2(n3201), .B1(n3491), .B2(
        \theRegs/completionDataOut[7][60] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[60].enDff/theFlop/N3 ) );
  AO22D0 U2933 ( .A1(n3555), .A2(n3200), .B1(n3635), .B2(
        \theRegs/completionDataOut[7][59] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[59].enDff/theFlop/N3 ) );
  AO22D0 U2934 ( .A1(n3436), .A2(n3199), .B1(n3498), .B2(
        \theRegs/completionDataOut[7][58] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[58].enDff/theFlop/N3 ) );
  AO22D0 U2935 ( .A1(n3764), .A2(n3198), .B1(n3809), .B2(
        \theRegs/completionDataOut[7][57] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[57].enDff/theFlop/N3 ) );
  AO22D0 U2937 ( .A1(n3555), .A2(n3179), .B1(n3392), .B2(
        \theRegs/completionDataOut[7][38] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[38].enDff/theFlop/N3 ) );
  AO22D0 U2938 ( .A1(n3572), .A2(n3178), .B1(n3652), .B2(
        \theRegs/completionDataOut[7][37] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[37].enDff/theFlop/N3 ) );
  AO22D0 U2939 ( .A1(n3862), .A2(n3177), .B1(n3911), .B2(
        \theRegs/completionDataOut[7][36] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[36].enDff/theFlop/N3 ) );
  AO22D0 U2940 ( .A1(n3566), .A2(n3194), .B1(n3685), .B2(
        \theRegs/completionDataOut[7][53] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[53].enDff/theFlop/N3 ) );
  AO22D0 U2941 ( .A1(n3764), .A2(n3193), .B1(n3809), .B2(
        \theRegs/completionDataOut[7][52] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[52].enDff/theFlop/N3 ) );
  AO22D0 U2943 ( .A1(n3536), .A2(n3192), .B1(n3735), .B2(
        \theRegs/completionDataOut[7][51] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[51].enDff/theFlop/N3 ) );
  AO22D0 U2944 ( .A1(n3566), .A2(n3191), .B1(n3685), .B2(
        \theRegs/completionDataOut[7][50] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[50].enDff/theFlop/N3 ) );
  AO22D0 U2945 ( .A1(n3989), .A2(n3190), .B1(n4017), .B2(
        \theRegs/completionDataOut[7][49] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[49].enDff/theFlop/N3 ) );
  AO22D0 U2946 ( .A1(n3632), .A2(n3189), .B1(n3777), .B2(
        \theRegs/completionDataOut[7][48] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[48].enDff/theFlop/N3 ) );
  AO22D0 U2947 ( .A1(n3566), .A2(n3188), .B1(n3504), .B2(
        \theRegs/completionDataOut[7][47] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[47].enDff/theFlop/N3 ) );
  AO22D0 U2948 ( .A1(n3860), .A2(n3187), .B1(n3910), .B2(
        \theRegs/completionDataOut[7][46] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[46].enDff/theFlop/N3 ) );
  AO22D0 U2949 ( .A1(n3722), .A2(n3186), .B1(n3775), .B2(
        \theRegs/completionDataOut[7][45] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[45].enDff/theFlop/N3 ) );
  AO22D0 U2950 ( .A1(n3436), .A2(n3185), .B1(n3635), .B2(
        \theRegs/completionDataOut[7][44] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[44].enDff/theFlop/N3 ) );
  AO22D0 U2951 ( .A1(n3555), .A2(n3184), .B1(n3635), .B2(
        \theRegs/completionDataOut[7][43] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[43].enDff/theFlop/N3 ) );
  AO22D0 U2952 ( .A1(n3722), .A2(n3183), .B1(n3775), .B2(
        \theRegs/completionDataOut[7][42] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[42].enDff/theFlop/N3 ) );
  AO22D0 U2953 ( .A1(n3425), .A2(n3182), .B1(n3491), .B2(
        \theRegs/completionDataOut[7][41] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[41].enDff/theFlop/N3 ) );
  AO22D0 U2954 ( .A1(n3740), .A2(n3181), .B1(n3797), .B2(
        \theRegs/completionDataOut[7][40] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[40].enDff/theFlop/N3 ) );
  AO22D0 U2955 ( .A1(n3376), .A2(n3180), .B1(n3392), .B2(
        \theRegs/completionDataOut[7][39] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[39].enDff/theFlop/N3 ) );
  AO22D0 U2957 ( .A1(n3572), .A2(n3146), .B1(n3652), .B2(
        \theRegs/completionDataOut[7][5] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U2958 ( .A1(n3572), .A2(n3145), .B1(n3652), .B2(
        \theRegs/completionDataOut[7][4] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U2959 ( .A1(n3740), .A2(n3144), .B1(n3797), .B2(
        \theRegs/completionDataOut[7][3] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U2960 ( .A1(n3722), .A2(n3176), .B1(n3498), .B2(
        \theRegs/completionDataOut[7][35] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[35].enDff/theFlop/N3 ) );
  AO22D0 U2961 ( .A1(n3376), .A2(n3175), .B1(n3491), .B2(
        \theRegs/completionDataOut[7][34] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[34].enDff/theFlop/N3 ) );
  AO22D0 U2963 ( .A1(n3632), .A2(n4045), .B1(n3777), .B2(
        \theRegs/completionDataOut[7][33] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[33].enDff/theFlop/N3 ) );
  AO22D0 U2964 ( .A1(n3566), .A2(n3173), .B1(n3504), .B2(
        \theRegs/completionDataOut[7][32] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[32].enDff/theFlop/N3 ) );
  AO22D0 U2965 ( .A1(n3566), .A2(n3172), .B1(n3504), .B2(
        \theRegs/completionDataOut[7][31] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[31].enDff/theFlop/N3 ) );
  AO22D0 U2966 ( .A1(n3632), .A2(n3171), .B1(n3504), .B2(
        \theRegs/completionDataOut[7][30] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[30].enDff/theFlop/N3 ) );
  AO22D0 U2967 ( .A1(n3860), .A2(n3170), .B1(n3910), .B2(
        \theRegs/completionDataOut[7][29] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[29].enDff/theFlop/N3 ) );
  AO22D0 U2968 ( .A1(n3602), .A2(n3169), .B1(n3777), .B2(
        \theRegs/completionDataOut[7][28] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[28].enDff/theFlop/N3 ) );
  AO22D0 U2969 ( .A1(n3764), .A2(n3168), .B1(n3809), .B2(
        \theRegs/completionDataOut[7][27] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[27].enDff/theFlop/N3 ) );
  AO22D0 U2970 ( .A1(n3903), .A2(n3167), .B1(n3952), .B2(
        \theRegs/completionDataOut[7][26] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[26].enDff/theFlop/N3 ) );
  AO22D0 U2971 ( .A1(n3903), .A2(n3166), .B1(n3952), .B2(
        \theRegs/completionDataOut[7][25] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[25].enDff/theFlop/N3 ) );
  AO22D0 U2972 ( .A1(n3903), .A2(n3165), .B1(n3952), .B2(
        \theRegs/completionDataOut[7][24] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[24].enDff/theFlop/N3 ) );
  AO22D0 U2973 ( .A1(n3764), .A2(n3164), .B1(n3809), .B2(
        \theRegs/completionDataOut[7][23] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[23].enDff/theFlop/N3 ) );
  AO22D0 U2974 ( .A1(n3989), .A2(n4092), .B1(n4017), .B2(
        \theRegs/completionDataOut[7][22] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[22].enDff/theFlop/N3 ) );
  AO22D0 U2975 ( .A1(n3566), .A2(n4112), .B1(n3504), .B2(
        \theRegs/completionDataOut[7][21] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[21].enDff/theFlop/N3 ) );
  AO22D0 U2976 ( .A1(n3989), .A2(n4113), .B1(n4017), .B2(
        \theRegs/completionDataOut[7][20] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[20].enDff/theFlop/N3 ) );
  AO22D0 U2977 ( .A1(n3331), .A2(n3160), .B1(n3316), .B2(
        \theRegs/completionDataOut[7][19] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[19].enDff/theFlop/N3 ) );
  AO22D0 U2978 ( .A1(n3632), .A2(n3159), .B1(n3504), .B2(
        \theRegs/completionDataOut[7][18] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[18].enDff/theFlop/N3 ) );
  AO22D0 U2980 ( .A1(n3536), .A2(n4048), .B1(n3735), .B2(
        \theRegs/completionDataOut[7][17] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[17].enDff/theFlop/N3 ) );
  AO22D0 U2981 ( .A1(n3903), .A2(n3157), .B1(n3952), .B2(
        \theRegs/completionDataOut[7][16] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[16].enDff/theFlop/N3 ) );
  AO22D0 U2984 ( .A1(n3764), .A2(n3156), .B1(n3809), .B2(
        \theRegs/completionDataOut[7][15] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[15].enDff/theFlop/N3 ) );
  AO22D0 U2985 ( .A1(n3989), .A2(n4054), .B1(n4017), .B2(
        \theRegs/completionDataOut[7][14] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[14].enDff/theFlop/N3 ) );
  AO22D0 U2986 ( .A1(n3860), .A2(n3154), .B1(n3910), .B2(
        \theRegs/completionDataOut[7][13] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[13].enDff/theFlop/N3 ) );
  AO22D0 U2987 ( .A1(n3764), .A2(n3153), .B1(n3809), .B2(
        \theRegs/completionDataOut[7][12] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[12].enDff/theFlop/N3 ) );
  AO22D0 U2988 ( .A1(n3602), .A2(n3152), .B1(n3777), .B2(
        \theRegs/completionDataOut[7][11] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[11].enDff/theFlop/N3 ) );
  AO22D0 U2989 ( .A1(n3536), .A2(n3151), .B1(n3735), .B2(
        \theRegs/completionDataOut[7][10] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[10].enDff/theFlop/N3 ) );
  AO22D0 U2990 ( .A1(n3632), .A2(n3150), .B1(n3777), .B2(
        \theRegs/completionDataOut[7][9] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[9].enDff/theFlop/N3 ) );
  AO22D0 U2991 ( .A1(n3602), .A2(n3149), .B1(n3735), .B2(
        \theRegs/completionDataOut[7][8] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U2992 ( .A1(n3860), .A2(n3148), .B1(n3910), .B2(
        \theRegs/completionDataOut[7][7] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U2993 ( .A1(n3903), .A2(n4089), .B1(n3952), .B2(
        \theRegs/completionDataOut[7][6] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U2994 ( .A1(n3862), .A2(n3142), .B1(n3911), .B2(
        \theRegs/completionDataOut[7][1] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U2995 ( .A1(n3740), .A2(n3143), .B1(n3797), .B2(
        \theRegs/completionDataOut[7][2] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U2996 ( .A1(n3436), .A2(n3141), .B1(n3498), .B2(
        \theRegs/completionDataOut[7][0] ), .Z(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U3006 ( .A1(n3223), .A2(n2211), .B1(n3690), .B2(
        \theRegs/managementDataOut[7][7] ), .Z(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U3007 ( .A1(n3221), .A2(n4039), .B1(n3762), .B2(
        \theRegs/managementDataOut[7][5] ), .Z(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U3008 ( .A1(n4043), .A2(n4039), .B1(n3762), .B2(
        \theRegs/managementDataOut[7][6] ), .Z(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U3009 ( .A1(n4096), .A2(n2211), .B1(n3690), .B2(
        \theRegs/managementDataOut[7][3] ), .Z(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U3010 ( .A1(n4042), .A2(n4039), .B1(n3690), .B2(
        \theRegs/managementDataOut[7][4] ), .Z(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U3011 ( .A1(n3986), .A2(n4039), .B1(n3762), .B2(
        \theRegs/managementDataOut[7][1] ), .Z(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U3012 ( .A1(n3900), .A2(n4039), .B1(n3762), .B2(
        \theRegs/managementDataOut[7][2] ), .Z(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U3013 ( .A1(n3901), .A2(n4039), .B1(n3762), .B2(
        \theRegs/managementDataOut[7][0] ), .Z(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U3019 ( .A1(n4096), .A2(n4033), .B1(n3753), .B2(
        \theRegs/managementDataOut[5][3] ), .Z(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U3020 ( .A1(n3900), .A2(n2219), .B1(n2218), .B2(
        \theRegs/managementDataOut[5][2] ), .Z(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U3021 ( .A1(n3986), .A2(n4033), .B1(n3753), .B2(
        \theRegs/managementDataOut[5][1] ), .Z(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U3022 ( .A1(n3216), .A2(n2219), .B1(n2218), .B2(
        \theRegs/managementDataOut[5][0] ), .Z(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U3023 ( .A1(n3899), .A2(n4033), .B1(n3753), .B2(
        \theRegs/managementDataOut[5][7] ), .Z(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U3024 ( .A1(n4043), .A2(n4033), .B1(n3753), .B2(
        \theRegs/managementDataOut[5][6] ), .Z(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U3025 ( .A1(n3221), .A2(n2219), .B1(n2218), .B2(
        \theRegs/managementDataOut[5][5] ), .Z(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U3026 ( .A1(n4042), .A2(n2219), .B1(n2218), .B2(
        \theRegs/managementDataOut[5][4] ), .Z(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U3027 ( .A1(n4012), .A2(n4033), .B1(\theRegs/managementDataOut[5][8] ), .B2(n3753), .Z(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U3030 ( .A1(n3220), .A2(n2226), .B1(n2225), .B2(
        \theRegs/managementDataOut[4][4] ), .Z(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U3031 ( .A1(n3222), .A2(n2226), .B1(n2225), .B2(
        \theRegs/managementDataOut[4][6] ), .Z(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U3032 ( .A1(n3899), .A2(n4032), .B1(n4116), .B2(
        \theRegs/managementDataOut[4][7] ), .Z(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U3033 ( .A1(n3901), .A2(n4032), .B1(n4116), .B2(
        \theRegs/managementDataOut[4][0] ), .Z(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U3034 ( .A1(n3902), .A2(n4032), .B1(n4116), .B2(
        \theRegs/managementDataOut[4][5] ), .Z(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U3035 ( .A1(n3900), .A2(n4032), .B1(n4116), .B2(
        \theRegs/managementDataOut[4][2] ), .Z(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U3036 ( .A1(n3219), .A2(n2226), .B1(n2225), .B2(
        \theRegs/managementDataOut[4][3] ), .Z(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U3037 ( .A1(n3986), .A2(n4032), .B1(n4116), .B2(
        \theRegs/managementDataOut[4][1] ), .Z(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U3038 ( .A1(n4012), .A2(n2226), .B1(\theRegs/managementDataOut[4][8] ), .B2(n4116), .Z(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U3042 ( .A1(n4013), .A2(\theRegs/managementDataOut[6][6] ), .B1(n3947), .B2(n3222), .Z(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U3043 ( .A1(n2215), .A2(\theRegs/managementDataOut[6][7] ), .B1(n2214), .B2(n3223), .Z(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U3044 ( .A1(n4013), .A2(\theRegs/managementDataOut[6][2] ), .B1(n3947), .B2(n3218), .Z(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U3045 ( .A1(n4013), .A2(\theRegs/managementDataOut[6][1] ), .B1(n2214), .B2(n3217), .Z(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U3046 ( .A1(n2215), .A2(\theRegs/managementDataOut[6][0] ), .B1(n2214), .B2(n3216), .Z(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U3047 ( .A1(n4013), .A2(\theRegs/managementDataOut[6][5] ), .B1(n2214), .B2(n3221), .Z(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U3048 ( .A1(n4013), .A2(\theRegs/managementDataOut[6][4] ), .B1(n3947), .B2(n3220), .Z(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U3049 ( .A1(n4013), .A2(\theRegs/managementDataOut[6][3] ), .B1(n3947), .B2(n3219), .Z(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U3050 ( .A1(\theRegs/managementDataOut[6][8] ), .A2(n2215), .B1(n3224), .B2(n3947), .Z(
        \theRegs/eachManagementReg[6].managementReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U3054 ( .A1(n4042), .A2(n2245), .B1(n3982), .B2(
        \theRegs/managementDataOut[0][4] ), .Z(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U3055 ( .A1(n3218), .A2(n2245), .B1(n3982), .B2(
        \theRegs/managementDataOut[0][2] ), .Z(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U3056 ( .A1(n3986), .A2(n4014), .B1(n4035), .B2(
        \theRegs/managementDataOut[0][1] ), .Z(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U3057 ( .A1(n3901), .A2(n2245), .B1(n3982), .B2(
        \theRegs/managementDataOut[0][0] ), .Z(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U3058 ( .A1(n4096), .A2(n4014), .B1(n4035), .B2(
        \theRegs/managementDataOut[0][3] ), .Z(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U3059 ( .A1(n3899), .A2(n4014), .B1(n4035), .B2(
        \theRegs/managementDataOut[0][7] ), .Z(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U3060 ( .A1(n4043), .A2(n4014), .B1(n4035), .B2(
        \theRegs/managementDataOut[0][6] ), .Z(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U3061 ( .A1(n3902), .A2(n4014), .B1(n4035), .B2(
        \theRegs/managementDataOut[0][5] ), .Z(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U3065 ( .A1(n3899), .A2(n2239), .B1(n2238), .B2(
        \theRegs/managementDataOut[1][7] ), .Z(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U3066 ( .A1(n4043), .A2(n4040), .B1(n2238), .B2(
        \theRegs/managementDataOut[1][6] ), .Z(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U3067 ( .A1(n4043), .A2(n3987), .B1(n3948), .B2(
        \theRegs/managementDataOut[2][6] ), .Z(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U3068 ( .A1(n3902), .A2(n3987), .B1(n3948), .B2(
        \theRegs/managementDataOut[2][5] ), .Z(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U3069 ( .A1(n3221), .A2(n2239), .B1(n2238), .B2(
        \theRegs/managementDataOut[1][5] ), .Z(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U3070 ( .A1(n4042), .A2(n4040), .B1(n4034), .B2(
        \theRegs/managementDataOut[1][4] ), .Z(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U3071 ( .A1(n4096), .A2(n2239), .B1(n2238), .B2(
        \theRegs/managementDataOut[1][3] ), .Z(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U3072 ( .A1(n3899), .A2(n3987), .B1(n2234), .B2(
        \theRegs/managementDataOut[2][7] ), .Z(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U3073 ( .A1(n3901), .A2(n3987), .B1(n3948), .B2(
        \theRegs/managementDataOut[2][0] ), .Z(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U3074 ( .A1(n3900), .A2(n4040), .B1(n4034), .B2(
        \theRegs/managementDataOut[1][2] ), .Z(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U3075 ( .A1(n3986), .A2(n4040), .B1(n4034), .B2(
        \theRegs/managementDataOut[1][1] ), .Z(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U3076 ( .A1(n3901), .A2(n4040), .B1(n4034), .B2(
        \theRegs/managementDataOut[1][0] ), .Z(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U3077 ( .A1(n4042), .A2(n3987), .B1(n3948), .B2(
        \theRegs/managementDataOut[2][4] ), .Z(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[4].enDff/theFlop/N3 ) );
  AO22D0 U3078 ( .A1(n4096), .A2(n2235), .B1(n2234), .B2(
        \theRegs/managementDataOut[2][3] ), .Z(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U3079 ( .A1(n3900), .A2(n2235), .B1(n2234), .B2(
        \theRegs/managementDataOut[2][2] ), .Z(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U3080 ( .A1(n3217), .A2(n2235), .B1(n2234), .B2(
        \theRegs/managementDataOut[2][1] ), .Z(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U3081 ( .A1(n4012), .A2(n2235), .B1(\theRegs/managementDataOut[2][8] ), .B2(n2234), .Z(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U3085 ( .A1(n4012), .A2(n2239), .B1(\theRegs/managementDataOut[1][8] ), .B2(n2238), .Z(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U3089 ( .A1(n4012), .A2(n2231), .B1(\theRegs/managementDataOut[3][8] ), .B2(n2230), .Z(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U3090 ( .A1(n3900), .A2(n3946), .B1(n3752), .B2(
        \theRegs/managementDataOut[3][2] ), .Z(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[2].enDff/theFlop/N3 ) );
  AO22D0 U3091 ( .A1(n3986), .A2(n3946), .B1(n3752), .B2(
        \theRegs/managementDataOut[3][1] ), .Z(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[1].enDff/theFlop/N3 ) );
  AO22D0 U3092 ( .A1(n3901), .A2(n3946), .B1(n3752), .B2(
        \theRegs/managementDataOut[3][0] ), .Z(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[0].enDff/theFlop/N3 ) );
  AO22D0 U3093 ( .A1(n4096), .A2(n2231), .B1(n2230), .B2(
        \theRegs/managementDataOut[3][3] ), .Z(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[3].enDff/theFlop/N3 ) );
  AO22D0 U3094 ( .A1(n3899), .A2(n2231), .B1(n2230), .B2(
        \theRegs/managementDataOut[3][7] ), .Z(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[7].enDff/theFlop/N3 ) );
  AO22D0 U3095 ( .A1(n4043), .A2(n3946), .B1(n3752), .B2(
        \theRegs/managementDataOut[3][6] ), .Z(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[6].enDff/theFlop/N3 ) );
  AO22D0 U3096 ( .A1(n3221), .A2(n2231), .B1(n2230), .B2(
        \theRegs/managementDataOut[3][5] ), .Z(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[5].enDff/theFlop/N3 ) );
  AO22D0 U3097 ( .A1(n4042), .A2(n3946), .B1(n3752), .B2(
        \theRegs/managementDataOut[3][4] ), .Z(
        \theRegs/eachManagementReg[3].managementReg/eachEnDff[4].enDff/theFlop/N3 ) );
  ND2D1 U4186 ( .A1(n3284), .A2(n3305), .ZN(n2246) );
  ND2D1 U4195 ( .A1(tail[0]), .A2(tail[1]), .ZN(n2203) );
  IND2D1 U4636 ( .A1(n2252), .B1(n2250), .ZN(n2257) );
  AO22D0 U4837 ( .A1(n4012), .A2(n2211), .B1(\theRegs/managementDataOut[7][8] ), .B2(n3690), .Z(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[8].enDff/theFlop/N3 ) );
  AO22D0 U4839 ( .A1(n3224), .A2(n2245), .B1(\theRegs/managementDataOut[0][8] ), .B2(n3982), .Z(
        \theRegs/eachManagementReg[0].managementReg/eachEnDff[8].enDff/theFlop/N3 ) );
  OA31D1 U4841 ( .A1(n3794), .A2(updateTail_i), .A3(
        \headTailManager/headReset ), .B(n2260), .Z(n1407) );
  NR2D1 U4842 ( .A1(n4031), .A2(n3794), .ZN(n2250) );
  AO211D1 U4845 ( .A1(n3247), .A2(n3874), .B(n4117), .C(n2252), .Z(n2253) );
  NR2XD1 U4175 ( .A1(n2224), .A2(n2223), .ZN(n2225) );
  NR3D8 U3018 ( .A1(n3242), .A2(n3246), .A3(n4041), .ZN(\add_x_7/n1 ) );
  MUX2ND1 U4836 ( .I0(tail[2]), .I1(n2265), .S(n2203), .ZN(n2207) );
  CKND2 U2660 ( .I(tail[0]), .ZN(n3238) );
  CKND12 U2662 ( .I(head[2]), .ZN(n3240) );
  BUFFD16 U2663 ( .I(head[1]), .Z(n3241) );
  CKND12 U2664 ( .I(n3241), .ZN(n3242) );
  BUFFD16 U2701 ( .I(head[0]), .Z(n3245) );
  CKND12 U2718 ( .I(n3245), .ZN(n3246) );
  BUFFD2 U2730 ( .I(head[0]), .Z(n3247) );
  CKND2 U2732 ( .I(n3247), .ZN(head_o[0]) );
  INVD1 U2783 ( .I(n3247), .ZN(n3250) );
  INVD1 U2962 ( .I(n2263), .ZN(n3283) );
  CKND3 U2979 ( .I(n3886), .ZN(n3284) );
  BUFFD16 U3064 ( .I(\add_x_7/n1 ), .Z(head_o[3]) );
  CKND3 U3087 ( .I(n3792), .ZN(n3306) );
  INVD1 U3088 ( .I(head_o[2]), .ZN(n3307) );
  ND4D8 U3481 ( .A1(n2442), .A2(n2441), .A3(n2440), .A4(n2439), .ZN(
        commitReadData_o[33]) );
  ND4D8 U3796 ( .A1(n2730), .A2(n2729), .A3(n2728), .A4(n2727), .ZN(
        decodeReadData1_o[32]) );
  ND4D8 U3786 ( .A1(n2722), .A2(n2721), .A3(n2720), .A4(n2719), .ZN(
        decodeReadData1_o[34]) );
  ND4D8 U3476 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), .ZN(
        commitReadData_o[34]) );
  ND4D8 U3951 ( .A1(n3003), .A2(n3002), .A3(n3001), .A4(n3000), .ZN(
        decodeReadData2_o[32]) );
  ND4D8 U3961 ( .A1(n2995), .A2(n2994), .A3(n2993), .A4(n2992), .ZN(
        decodeReadData2_o[34]) );
  ND4D8 U3486 ( .A1(n2438), .A2(n2437), .A3(n2436), .A4(n2435), .ZN(
        commitReadData_o[32]) );
  ND4D8 U3791 ( .A1(n2726), .A2(n2725), .A3(n2724), .A4(n2723), .ZN(
        decodeReadData1_o[33]) );
  ND4D8 U3956 ( .A1(n2999), .A2(n2998), .A3(n2997), .A4(n2996), .ZN(
        decodeReadData2_o[33]) );
  ND4D8 U3441 ( .A1(n2474), .A2(n2473), .A3(n2472), .A4(n2471), .ZN(
        commitReadData_o[41]) );
  ND4D8 U3491 ( .A1(n2434), .A2(n2433), .A3(n2432), .A4(n2431), .ZN(
        commitReadData_o[31]) );
  ND4D8 U3946 ( .A1(n3007), .A2(n3006), .A3(n3005), .A4(n3004), .ZN(
        decodeReadData2_o[31]) );
  ND4D8 U3801 ( .A1(n2734), .A2(n2733), .A3(n2732), .A4(n2731), .ZN(
        decodeReadData1_o[31]) );
  ND4D8 U3496 ( .A1(n2430), .A2(n2429), .A3(n2428), .A4(n2427), .ZN(
        commitReadData_o[30]) );
  ND4D8 U3941 ( .A1(n3011), .A2(n3010), .A3(n3009), .A4(n3008), .ZN(
        decodeReadData2_o[30]) );
  ND4D8 U3966 ( .A1(n2991), .A2(n2990), .A3(n2989), .A4(n2988), .ZN(
        decodeReadData2_o[35]) );
  ND4D8 U3806 ( .A1(n2738), .A2(n2737), .A3(n2736), .A4(n2735), .ZN(
        decodeReadData1_o[30]) );
  ND4D8 U3781 ( .A1(n2718), .A2(n2717), .A3(n2716), .A4(n2715), .ZN(
        decodeReadData1_o[35]) );
  ND4D8 U3816 ( .A1(n2746), .A2(n2745), .A3(n2744), .A4(n2743), .ZN(
        decodeReadData1_o[28]) );
  ND4D8 U4006 ( .A1(n3015), .A2(n3014), .A3(n3013), .A4(n3012), .ZN(
        decodeReadData2_o[29]) );
  ND4D8 U3501 ( .A1(n2426), .A2(n2425), .A3(n2424), .A4(n2423), .ZN(
        commitReadData_o[29]) );
  ND4D8 U3701 ( .A1(n2658), .A2(n2657), .A3(n2656), .A4(n2655), .ZN(
        decodeReadData1_o[50]) );
  ND4D8 U3446 ( .A1(n2470), .A2(n2469), .A3(n2468), .A4(n2467), .ZN(
        commitReadData_o[40]) );
  ND4D8 U3811 ( .A1(n2742), .A2(n2741), .A3(n2740), .A4(n2739), .ZN(
        decodeReadData1_o[29]) );
  ND4D8 U3506 ( .A1(n2422), .A2(n2421), .A3(n2420), .A4(n2419), .ZN(
        commitReadData_o[28]) );
  ND4D8 U3401 ( .A1(n2506), .A2(n2505), .A3(n2504), .A4(n2503), .ZN(
        commitReadData_o[49]) );
  ND4D8 U3356 ( .A1(n3019), .A2(n3018), .A3(n3017), .A4(n3016), .ZN(
        decodeReadData2_o[28]) );
  ND4D8 U3396 ( .A1(n2510), .A2(n2509), .A3(n2508), .A4(n2507), .ZN(
        commitReadData_o[50]) );
  ND4D8 U4046 ( .A1(n2931), .A2(n2930), .A3(n2929), .A4(n2928), .ZN(
        decodeReadData2_o[50]) );
  ND4D8 U3651 ( .A1(n2666), .A2(n2665), .A3(n2664), .A4(n2663), .ZN(
        decodeReadData1_o[48]) );
  ND4D8 U3996 ( .A1(n2971), .A2(n2970), .A3(n2969), .A4(n2968), .ZN(
        decodeReadData2_o[40]) );
  ND4D8 U3691 ( .A1(n2698), .A2(n2697), .A3(n2696), .A4(n2695), .ZN(
        decodeReadData1_o[40]) );
  ND4D8 U4041 ( .A1(n2935), .A2(n2934), .A3(n2933), .A4(n2932), .ZN(
        decodeReadData2_o[49]) );
  ND4D8 U4036 ( .A1(n2939), .A2(n2938), .A3(n2937), .A4(n2936), .ZN(
        decodeReadData2_o[48]) );
  ND4D8 U3661 ( .A1(n2674), .A2(n2673), .A3(n2672), .A4(n2671), .ZN(
        decodeReadData1_o[46]) );
  ND4D8 U3416 ( .A1(n2494), .A2(n2493), .A3(n2492), .A4(n2491), .ZN(
        commitReadData_o[46]) );
  ND4D8 U4026 ( .A1(n2947), .A2(n2946), .A3(n2945), .A4(n2944), .ZN(
        decodeReadData2_o[46]) );
  ND4D8 U3686 ( .A1(n2694), .A2(n2693), .A3(n2692), .A4(n2691), .ZN(
        decodeReadData1_o[41]) );
  ND4D8 U3681 ( .A1(n2690), .A2(n2689), .A3(n2688), .A4(n2687), .ZN(
        decodeReadData1_o[42]) );
  ND4D8 U3751 ( .A1(n2662), .A2(n2661), .A3(n2660), .A4(n2659), .ZN(
        decodeReadData1_o[49]) );
  ND4D8 U4031 ( .A1(n2943), .A2(n2942), .A3(n2941), .A4(n2940), .ZN(
        decodeReadData2_o[47]) );
  ND4D8 U3656 ( .A1(n2670), .A2(n2669), .A3(n2668), .A4(n2667), .ZN(
        decodeReadData1_o[47]) );
  ND4D8 U4021 ( .A1(n2951), .A2(n2950), .A3(n2949), .A4(n2948), .ZN(
        decodeReadData2_o[45]) );
  ND4D8 U4001 ( .A1(n2967), .A2(n2966), .A3(n2965), .A4(n2964), .ZN(
        decodeReadData2_o[41]) );
  ND4D8 U3511 ( .A1(n2418), .A2(n2417), .A3(n2416), .A4(n2415), .ZN(
        commitReadData_o[27]) );
  ND4D8 U4086 ( .A1(n2963), .A2(n2962), .A3(n2961), .A4(n2960), .ZN(
        decodeReadData2_o[42]) );
  ND4D8 U3711 ( .A1(n2650), .A2(n2649), .A3(n2648), .A4(n2647), .ZN(
        decodeReadData1_o[52]) );
  ND4D8 U3406 ( .A1(n2502), .A2(n2501), .A3(n2500), .A4(n2499), .ZN(
        commitReadData_o[48]) );
  ND4D8 U3821 ( .A1(n2750), .A2(n2749), .A3(n2748), .A4(n2747), .ZN(
        decodeReadData1_o[27]) );
  ND4D8 U3110 ( .A1(n3023), .A2(n3022), .A3(n3021), .A4(n3020), .ZN(
        decodeReadData2_o[27]) );
  ND4D8 U3706 ( .A1(n2654), .A2(n2653), .A3(n2652), .A4(n2651), .ZN(
        decodeReadData1_o[51]) );
  ND4D8 U3411 ( .A1(n2498), .A2(n2497), .A3(n2496), .A4(n2495), .ZN(
        commitReadData_o[47]) );
  ND4D8 U3436 ( .A1(n2478), .A2(n2477), .A3(n2476), .A4(n2475), .ZN(
        commitReadData_o[42]) );
  ND4D8 U3431 ( .A1(n2482), .A2(n2481), .A3(n2480), .A4(n2479), .ZN(
        commitReadData_o[43]) );
  ND4D8 U3676 ( .A1(n2686), .A2(n2685), .A3(n2684), .A4(n2683), .ZN(
        decodeReadData1_o[43]) );
  ND4D8 U3826 ( .A1(n2754), .A2(n2753), .A3(n2752), .A4(n2751), .ZN(
        decodeReadData1_o[26]) );
  ND4D8 U4101 ( .A1(n2866), .A2(n2865), .A3(n2864), .A4(n2863), .ZN(
        decodeReadData1_o[0]) );
  ND4D8 U3666 ( .A1(n2678), .A2(n2677), .A3(n2676), .A4(n2675), .ZN(
        decodeReadData1_o[45]) );
  ND4D8 U3766 ( .A1(n2706), .A2(n2705), .A3(n2704), .A4(n2703), .ZN(
        decodeReadData1_o[38]) );
  ND4D8 U3386 ( .A1(n2518), .A2(n2517), .A3(n2516), .A4(n2515), .ZN(
        commitReadData_o[52]) );
  ND4D8 U4056 ( .A1(n2923), .A2(n2922), .A3(n2921), .A4(n2920), .ZN(
        decodeReadData2_o[52]) );
  ND4D8 U3421 ( .A1(n2490), .A2(n2489), .A3(n2488), .A4(n2487), .ZN(
        commitReadData_o[45]) );
  ND4D8 U3115 ( .A1(n3027), .A2(n3026), .A3(n3025), .A4(n3024), .ZN(
        decodeReadData2_o[26]) );
  ND4D8 U3426 ( .A1(n2486), .A2(n2485), .A3(n2484), .A4(n2483), .ZN(
        commitReadData_o[44]) );
  ND4D8 U4051 ( .A1(n2927), .A2(n2926), .A3(n2925), .A4(n2924), .ZN(
        decodeReadData2_o[51]) );
  ND4D8 U3671 ( .A1(n2682), .A2(n2681), .A3(n2680), .A4(n2679), .ZN(
        decodeReadData1_o[44]) );
  ND4D8 U4016 ( .A1(n2955), .A2(n2954), .A3(n2953), .A4(n2952), .ZN(
        decodeReadData2_o[44]) );
  ND4D8 U4011 ( .A1(n2959), .A2(n2958), .A3(n2957), .A4(n2956), .ZN(
        decodeReadData2_o[43]) );
  ND4D8 U3831 ( .A1(n2758), .A2(n2757), .A3(n2756), .A4(n2755), .ZN(
        decodeReadData1_o[25]) );
  ND4D8 U3696 ( .A1(n2702), .A2(n2701), .A3(n2700), .A4(n2699), .ZN(
        decodeReadData1_o[39]) );
  ND4D8 U3120 ( .A1(n3031), .A2(n3030), .A3(n3029), .A4(n3028), .ZN(
        decodeReadData2_o[25]) );
  ND4D8 U3516 ( .A1(n2414), .A2(n2413), .A3(n2412), .A4(n2411), .ZN(
        commitReadData_o[26]) );
  ND4D8 U3391 ( .A1(n2514), .A2(n2513), .A3(n2512), .A4(n2511), .ZN(
        commitReadData_o[51]) );
  ND4D8 U3771 ( .A1(n2710), .A2(n2709), .A3(n2708), .A4(n2707), .ZN(
        decodeReadData1_o[37]) );
  ND4D8 U3986 ( .A1(n2979), .A2(n2978), .A3(n2977), .A4(n2976), .ZN(
        decodeReadData2_o[38]) );
  ND4D8 U3776 ( .A1(n2714), .A2(n2713), .A3(n2712), .A4(n2711), .ZN(
        decodeReadData1_o[36]) );
  NR2D3 U4826 ( .A1(n2236), .A2(n2237), .ZN(n2239) );
  ND4D8 U3381 ( .A1(n2522), .A2(n2521), .A3(n2520), .A4(n2519), .ZN(
        commitReadData_o[53]) );
  ND4D8 U3601 ( .A1(n2346), .A2(n2345), .A3(n2344), .A4(n2343), .ZN(
        commitReadData_o[9]) );
  ND4D8 U3606 ( .A1(n2342), .A2(n2341), .A3(n2340), .A4(n2339), .ZN(
        commitReadData_o[8]) );
  ND4D8 U3521 ( .A1(n2410), .A2(n2409), .A3(n2408), .A4(n2407), .ZN(
        commitReadData_o[25]) );
  ND4D8 U3245 ( .A1(n3139), .A2(n3138), .A3(n3137), .A4(n3136), .ZN(
        decodeReadData2_o[0]) );
  ND4D8 U3581 ( .A1(n2362), .A2(n2361), .A3(n2360), .A4(n2359), .ZN(
        commitReadData_o[13]) );
  ND4D8 U3576 ( .A1(n2366), .A2(n2365), .A3(n2364), .A4(n2363), .ZN(
        commitReadData_o[14]) );
  ND4D8 U3596 ( .A1(n2350), .A2(n2349), .A3(n2348), .A4(n2347), .ZN(
        commitReadData_o[10]) );
  ND4D8 U3125 ( .A1(n3035), .A2(n3034), .A3(n3033), .A4(n3032), .ZN(
        decodeReadData2_o[24]) );
  ND4D8 U3616 ( .A1(n2334), .A2(n2333), .A3(n2332), .A4(n2331), .ZN(
        commitReadData_o[6]) );
  ND4D8 U3841 ( .A1(n2766), .A2(n2765), .A3(n2764), .A4(n2763), .ZN(
        decodeReadData1_o[23]) );
  ND4D8 U3571 ( .A1(n2370), .A2(n2369), .A3(n2368), .A4(n2367), .ZN(
        commitReadData_o[15]) );
  ND4D8 U3976 ( .A1(n2983), .A2(n2982), .A3(n2981), .A4(n2980), .ZN(
        decodeReadData2_o[37]) );
  ND4D8 U3971 ( .A1(n2987), .A2(n2986), .A3(n2985), .A4(n2984), .ZN(
        decodeReadData2_o[36]) );
  ND4D8 U3240 ( .A1(n3127), .A2(n3126), .A3(n3125), .A4(n3124), .ZN(
        decodeReadData2_o[1]) );
  ND4D8 U3230 ( .A1(n3119), .A2(n3118), .A3(n3117), .A4(n3116), .ZN(
        decodeReadData2_o[3]) );
  ND4D8 U3180 ( .A1(n3079), .A2(n3078), .A3(n3077), .A4(n3076), .ZN(
        decodeReadData2_o[13]) );
  ND4D8 U3195 ( .A1(n3091), .A2(n3090), .A3(n3089), .A4(n3088), .ZN(
        decodeReadData2_o[10]) );
  ND4D8 U3210 ( .A1(n3103), .A2(n3102), .A3(n3101), .A4(n3100), .ZN(
        decodeReadData2_o[7]) );
  ND4D8 U3836 ( .A1(n2762), .A2(n2761), .A3(n2760), .A4(n2759), .ZN(
        decodeReadData1_o[24]) );
  ND4D8 U3205 ( .A1(n3099), .A2(n3098), .A3(n3097), .A4(n3096), .ZN(
        decodeReadData2_o[8]) );
  ND4D8 U3586 ( .A1(n2358), .A2(n2357), .A3(n2356), .A4(n2355), .ZN(
        commitReadData_o[12]) );
  ND4D8 U3200 ( .A1(n3095), .A2(n3094), .A3(n3093), .A4(n3092), .ZN(
        decodeReadData2_o[9]) );
  ND4D8 U3130 ( .A1(n3039), .A2(n3038), .A3(n3037), .A4(n3036), .ZN(
        decodeReadData2_o[23]) );
  ND4D8 U3185 ( .A1(n3083), .A2(n3082), .A3(n3081), .A4(n3080), .ZN(
        decodeReadData2_o[12]) );
  ND4D8 U4061 ( .A1(n2919), .A2(n2918), .A3(n2917), .A4(n2916), .ZN(
        decodeReadData2_o[53]) );
  ND4D8 U3991 ( .A1(n2975), .A2(n2974), .A3(n2973), .A4(n2972), .ZN(
        decodeReadData2_o[39]) );
  ND4D8 U3916 ( .A1(n2826), .A2(n2825), .A3(n2824), .A4(n2823), .ZN(
        decodeReadData1_o[8]) );
  NR2D3 U4182 ( .A1(n2240), .A2(n2241), .ZN(n2245) );
  ND4D8 U3896 ( .A1(n2810), .A2(n2809), .A3(n2808), .A4(n2807), .ZN(
        decodeReadData1_o[12]) );
  ND4D8 U3561 ( .A1(n2378), .A2(n2377), .A3(n2376), .A4(n2375), .ZN(
        commitReadData_o[17]) );
  ND4D8 U3321 ( .A1(n2566), .A2(n2565), .A3(n2564), .A4(n2563), .ZN(
        commitReadData_o[64]) );
  ND4D8 U3225 ( .A1(n3115), .A2(n3114), .A3(n3113), .A4(n3112), .ZN(
        decodeReadData2_o[4]) );
  ND4D8 U3906 ( .A1(n2818), .A2(n2817), .A3(n2816), .A4(n2815), .ZN(
        decodeReadData1_o[10]) );
  ND4D8 U3921 ( .A1(n2830), .A2(n2829), .A3(n2828), .A4(n2827), .ZN(
        decodeReadData1_o[7]) );
  ND4D8 U3531 ( .A1(n2402), .A2(n2401), .A3(n2400), .A4(n2399), .ZN(
        commitReadData_o[23]) );
  ND4D8 U3911 ( .A1(n2822), .A2(n2821), .A3(n2820), .A4(n2819), .ZN(
        decodeReadData1_o[9]) );
  ND4D8 U3215 ( .A1(n3107), .A2(n3106), .A3(n3105), .A4(n3104), .ZN(
        decodeReadData2_o[6]) );
  ND4D8 U4121 ( .A1(n2618), .A2(n2617), .A3(n2616), .A4(n2615), .ZN(
        decodeReadData1_o[60]) );
  ND4D8 U3376 ( .A1(n2526), .A2(n2525), .A3(n2524), .A4(n2523), .ZN(
        commitReadData_o[54]) );
  ND4D8 U4106 ( .A1(n2854), .A2(n2853), .A3(n2852), .A4(n2851), .ZN(
        decodeReadData1_o[1]) );
  ND4D8 U3220 ( .A1(n3111), .A2(n3110), .A3(n3109), .A4(n3108), .ZN(
        decodeReadData2_o[5]) );
  ND4D8 U3566 ( .A1(n2374), .A2(n2373), .A3(n2372), .A4(n2371), .ZN(
        commitReadData_o[16]) );
  ND4D8 U4116 ( .A1(n2846), .A2(n2845), .A3(n2844), .A4(n2843), .ZN(
        decodeReadData1_o[3]) );
  ND4D8 U3235 ( .A1(n3123), .A2(n3122), .A3(n3121), .A4(n3120), .ZN(
        decodeReadData2_o[2]) );
  DFQD4 \headTailManager/head_reg[2]  ( .D(n1404), .CP(clk_i), .Q(head[2]) );
  ND4D8 U3526 ( .A1(n2406), .A2(n2405), .A3(n2404), .A4(n2403), .ZN(
        commitReadData_o[24]) );
  ND4D8 U3716 ( .A1(n2646), .A2(n2645), .A3(n2644), .A4(n2643), .ZN(
        decodeReadData1_o[53]) );
  ND4D8 U3891 ( .A1(n2806), .A2(n2805), .A3(n2804), .A4(n2803), .ZN(
        decodeReadData1_o[13]) );
  ND4D8 U3165 ( .A1(n3067), .A2(n3066), .A3(n3065), .A4(n3064), .ZN(
        decodeReadData2_o[16]) );
  ND4D8 U4096 ( .A1(n2875), .A2(n2874), .A3(n2873), .A4(n2872), .ZN(
        decodeReadData2_o[64]) );
  ND4D8 U3170 ( .A1(n3071), .A2(n3070), .A3(n3069), .A4(n3068), .ZN(
        decodeReadData2_o[15]) );
  ND4D8 U3591 ( .A1(n2354), .A2(n2353), .A3(n2352), .A4(n2351), .ZN(
        commitReadData_o[11]) );
  ND4D8 U3336 ( .A1(n2554), .A2(n2553), .A3(n2552), .A4(n2551), .ZN(
        commitReadData_o[61]) );
  ND4D8 U3931 ( .A1(n2838), .A2(n2837), .A3(n2836), .A4(n2835), .ZN(
        decodeReadData1_o[5]) );
  NR3D8 U4177 ( .A1(n3240), .A2(n3241), .A3(n3245), .ZN(n2583) );
  ND4D8 U3160 ( .A1(n3063), .A2(n3062), .A3(n3061), .A4(n3060), .ZN(
        decodeReadData2_o[17]) );
  ND4D8 U3926 ( .A1(n2834), .A2(n2833), .A3(n2832), .A4(n2831), .ZN(
        decodeReadData1_o[6]) );
  ND4D8 U3536 ( .A1(n2398), .A2(n2397), .A3(n2396), .A4(n2395), .ZN(
        commitReadData_o[22]) );
  ND4D8 U3190 ( .A1(n3087), .A2(n3086), .A3(n3085), .A4(n3084), .ZN(
        decodeReadData2_o[11]) );
  ND4D8 U4139 ( .A1(n2891), .A2(n2890), .A3(n2889), .A4(n2888), .ZN(
        decodeReadData2_o[60]) );
  ND4D8 U4111 ( .A1(n2850), .A2(n2849), .A3(n2848), .A4(n2847), .ZN(
        decodeReadData1_o[2]) );
  ND4D8 U3175 ( .A1(n3075), .A2(n3074), .A3(n3073), .A4(n3072), .ZN(
        decodeReadData2_o[14]) );
  ND4D8 U3981 ( .A1(n2602), .A2(n2601), .A3(n2600), .A4(n2599), .ZN(
        decodeReadData1_o[64]) );
  ND4D8 U3871 ( .A1(n2790), .A2(n2789), .A3(n2788), .A4(n2787), .ZN(
        decodeReadData1_o[17]) );
  ND4D8 U3936 ( .A1(n2842), .A2(n2841), .A3(n2840), .A4(n2839), .ZN(
        decodeReadData1_o[4]) );
  ND4D8 U4066 ( .A1(n2915), .A2(n2914), .A3(n2913), .A4(n2912), .ZN(
        decodeReadData2_o[54]) );
  ND4D8 U3556 ( .A1(n2382), .A2(n2381), .A3(n2380), .A4(n2379), .ZN(
        commitReadData_o[18]) );
  ND4D8 U3881 ( .A1(n2798), .A2(n2797), .A3(n2796), .A4(n2795), .ZN(
        decodeReadData1_o[15]) );
  ND4D8 U3846 ( .A1(n2770), .A2(n2769), .A3(n2768), .A4(n2767), .ZN(
        decodeReadData1_o[22]) );
  ND4D8 U3876 ( .A1(n2794), .A2(n2793), .A3(n2792), .A4(n2791), .ZN(
        decodeReadData1_o[16]) );
  ND4D8 U3351 ( .A1(n2542), .A2(n2541), .A3(n2540), .A4(n2539), .ZN(
        commitReadData_o[58]) );
  ND4D8 U3901 ( .A1(n2814), .A2(n2813), .A3(n2812), .A4(n2811), .ZN(
        decodeReadData1_o[11]) );
  ND4D8 U3721 ( .A1(n2642), .A2(n2641), .A3(n2640), .A4(n2639), .ZN(
        decodeReadData1_o[54]) );
  ND4D8 U3341 ( .A1(n2550), .A2(n2549), .A3(n2548), .A4(n2547), .ZN(
        commitReadData_o[60]) );
  ND4D8 U3366 ( .A1(n2534), .A2(n2533), .A3(n2532), .A4(n2531), .ZN(
        commitReadData_o[56]) );
  ND4D8 U3155 ( .A1(n3059), .A2(n3058), .A3(n3057), .A4(n3056), .ZN(
        decodeReadData2_o[18]) );
  ND4D8 U3326 ( .A1(n2562), .A2(n2561), .A3(n2560), .A4(n2559), .ZN(
        commitReadData_o[63]) );
  ND4D8 U3756 ( .A1(n2614), .A2(n2613), .A3(n2612), .A4(n2611), .ZN(
        decodeReadData1_o[61]) );
  ND4D8 U3646 ( .A1(n2606), .A2(n2605), .A3(n2604), .A4(n2603), .ZN(
        decodeReadData1_o[63]) );
  ND4D8 U3886 ( .A1(n2802), .A2(n2801), .A3(n2800), .A4(n2799), .ZN(
        decodeReadData1_o[14]) );
  ND4D8 U3331 ( .A1(n2558), .A2(n2557), .A3(n2556), .A4(n2555), .ZN(
        commitReadData_o[62]) );
  ND4D8 U3866 ( .A1(n2786), .A2(n2785), .A3(n2784), .A4(n2783), .ZN(
        decodeReadData1_o[18]) );
  INR2XD1 U4256 ( .A1(n2270), .B1(n3974), .ZN(stall_o) );
  ND4D8 U4144 ( .A1(n2887), .A2(n2886), .A3(n2885), .A4(n2884), .ZN(
        decodeReadData2_o[61]) );
  ND4D8 U3551 ( .A1(n2386), .A2(n2385), .A3(n2384), .A4(n2383), .ZN(
        commitReadData_o[19]) );
  ND4D8 U4149 ( .A1(n2895), .A2(n2894), .A3(n2893), .A4(n2892), .ZN(
        decodeReadData2_o[59]) );
  ND4D8 U3746 ( .A1(n2622), .A2(n2621), .A3(n2620), .A4(n2619), .ZN(
        decodeReadData1_o[59]) );
  ND4D8 U3541 ( .A1(n2394), .A2(n2393), .A3(n2392), .A4(n2391), .ZN(
        commitReadData_o[21]) );
  ND4D8 U3361 ( .A1(n2538), .A2(n2537), .A3(n2536), .A4(n2535), .ZN(
        commitReadData_o[57]) );
  ND4D8 U3135 ( .A1(n3043), .A2(n3042), .A3(n3041), .A4(n3040), .ZN(
        decodeReadData2_o[22]) );
  BUFFD2 U2289 ( .I(completionWriteData_i[18]), .Z(n3159) );
  ND4D8 U3371 ( .A1(n2530), .A2(n2529), .A3(n2528), .A4(n2527), .ZN(
        commitReadData_o[55]) );
  ND4D8 U3731 ( .A1(n2634), .A2(n2633), .A3(n2632), .A4(n2631), .ZN(
        decodeReadData1_o[56]) );
  BUFFD2 U2291 ( .I(completionWriteData_i[20]), .Z(n3161) );
  BUFFD2 U2292 ( .I(completionWriteData_i[21]), .Z(n3162) );
  ND4D8 U4091 ( .A1(n2899), .A2(n2898), .A3(n2897), .A4(n2896), .ZN(
        decodeReadData2_o[58]) );
  ND4D8 U3546 ( .A1(n2390), .A2(n2389), .A3(n2388), .A4(n2387), .ZN(
        commitReadData_o[20]) );
  ND4D8 U3726 ( .A1(n2638), .A2(n2637), .A3(n2636), .A4(n2635), .ZN(
        decodeReadData1_o[55]) );
  ND4D8 U3761 ( .A1(n2610), .A2(n2609), .A3(n2608), .A4(n2607), .ZN(
        decodeReadData1_o[62]) );
  ND4D8 U4134 ( .A1(n2879), .A2(n2878), .A3(n2877), .A4(n2876), .ZN(
        decodeReadData2_o[63]) );
  ND4D8 U4081 ( .A1(n2903), .A2(n2902), .A3(n2901), .A4(n2900), .ZN(
        decodeReadData2_o[57]) );
  ND4D8 U3736 ( .A1(n2630), .A2(n2629), .A3(n2628), .A4(n2627), .ZN(
        decodeReadData1_o[57]) );
  ND4D8 U4071 ( .A1(n2911), .A2(n2910), .A3(n2909), .A4(n2908), .ZN(
        decodeReadData2_o[55]) );
  NR2D1 U4197 ( .A1(n3227), .A2(n2871), .ZN(n3134) );
  ND4D8 U3346 ( .A1(n2546), .A2(n2545), .A3(n2544), .A4(n2543), .ZN(
        commitReadData_o[59]) );
  ND4D2 U3741 ( .A1(n2626), .A2(n2625), .A3(n2624), .A4(n2623), .ZN(
        decodeReadData1_o[58]) );
  ND4D8 U4076 ( .A1(n2907), .A2(n2906), .A3(n2905), .A4(n2904), .ZN(
        decodeReadData2_o[56]) );
  ND4D8 U3150 ( .A1(n3055), .A2(n3054), .A3(n3053), .A4(n3052), .ZN(
        decodeReadData2_o[19]) );
  AOI22D2 U3262 ( .A1(n3297), .A2(\theRegs/managementDataOut[6][6] ), .B1(
        head_o[3]), .B2(\theRegs/managementDataOut[7][6] ), .ZN(n2295) );
  BUFFD2 U2297 ( .I(completionWriteData_i[25]), .Z(n3166) );
  BUFFD2 U2299 ( .I(completionWriteData_i[26]), .Z(n3167) );
  ND4D8 U4129 ( .A1(n2883), .A2(n2882), .A3(n2881), .A4(n2880), .ZN(
        decodeReadData2_o[62]) );
  BUFFD2 U2300 ( .I(completionWriteData_i[27]), .Z(n3168) );
  BUFFD2 U2322 ( .I(completionWriteData_i[44]), .Z(n3185) );
  BUFFD2 U2325 ( .I(completionWriteData_i[47]), .Z(n3188) );
  BUFFD2 U2310 ( .I(completionWriteData_i[35]), .Z(n3176) );
  BUFFD2 U2302 ( .I(completionWriteData_i[29]), .Z(n3170) );
  BUFFD2 U2308 ( .I(completionWriteData_i[34]), .Z(n3175) );
  AOI22D2 U3265 ( .A1(n3300), .A2(\theRegs/managementDataOut[5][6] ), .B1(
        n3298), .B2(\theRegs/managementDataOut[4][6] ), .ZN(n2298) );
  ND4D8 U3145 ( .A1(n3051), .A2(n3050), .A3(n3049), .A4(n3048), .ZN(
        decodeReadData2_o[20]) );
  BUFFD2 U2301 ( .I(completionWriteData_i[28]), .Z(n3169) );
  BUFFD2 U2327 ( .I(completionWriteData_i[49]), .Z(n3190) );
  BUFFD2 U2318 ( .I(completionWriteData_i[40]), .Z(n3181) );
  BUFFD2 U2321 ( .I(completionWriteData_i[43]), .Z(n3184) );
  NR2D4 U4820 ( .A1(n2208), .A2(n3885), .ZN(n2211) );
  BUFFD2 U2276 ( .I(completionWriteData_i[11]), .Z(n3152) );
  BUFFD1 U2296 ( .I(completionWriteData_i[24]), .Z(n3165) );
  BUFFD2 U2319 ( .I(completionWriteData_i[41]), .Z(n3182) );
  BUFFD1 U2498 ( .I(decodeWriteData_i[3]), .Z(n3219) );
  BUFFD2 U2320 ( .I(completionWriteData_i[42]), .Z(n3183) );
  BUFFD2 U2323 ( .I(completionWriteData_i[45]), .Z(n3186) );
  BUFFD2 U2295 ( .I(completionWriteData_i[23]), .Z(n3164) );
  BUFFD2 U2294 ( .I(completionWriteData_i[22]), .Z(n3163) );
  BUFFD2 U2274 ( .I(completionWriteData_i[10]), .Z(n3151) );
  INR2XD2 U3086 ( .A1(n2237), .B1(n2236), .ZN(n2238) );
  AOI22D2 U3300 ( .A1(n3300), .A2(\theRegs/completionDataOut[5][69] ), .B1(
        n3298), .B2(\theRegs/completionDataOut[4][69] ), .ZN(n2593) );
  BUFFD2 U2269 ( .I(completionWriteData_i[7]), .Z(n3148) );
  BUFFD2 U2268 ( .I(completionWriteData_i[6]), .Z(n3147) );
  BUFFD2 U2264 ( .I(completionWriteData_i[3]), .Z(n3144) );
  BUFFD2 U2273 ( .I(completionWriteData_i[9]), .Z(n3150) );
  BUFFD2 U2393 ( .I(completionWriteData_i[57]), .Z(n3198) );
  AOI22D2 U3632 ( .A1(n3297), .A2(\theRegs/completionDataOut[6][3] ), .B1(
        head_o[3]), .B2(\theRegs/completionDataOut[7][3] ), .ZN(n2319) );
  BUFFD2 U2332 ( .I(completionWriteData_i[54]), .Z(n3195) );
  BUFFD2 U2271 ( .I(completionWriteData_i[8]), .Z(n3149) );
  BUFFD2 U2262 ( .I(completionWriteData_i[1]), .Z(n3142) );
  BUFFD2 U2392 ( .I(completionWriteData_i[56]), .Z(n3197) );
  BUFFD1 U2316 ( .I(completionWriteData_i[39]), .Z(n3180) );
  AOI22D2 U3252 ( .A1(\theRegs/managementDataOut[6][8] ), .A2(n3297), .B1(
        \theRegs/managementDataOut[7][8] ), .B2(n3703), .ZN(n2303) );
  BUFFD2 U2265 ( .I(completionWriteData_i[4]), .Z(n3145) );
  BUFFD2 U2263 ( .I(completionWriteData_i[2]), .Z(n3143) );
  BUFFD2 U2407 ( .I(completionWriteData_i[60]), .Z(n3201) );
  BUFFD1 U2313 ( .I(completionWriteData_i[37]), .Z(n3178) );
  BUFFD2 U2324 ( .I(completionWriteData_i[46]), .Z(n3187) );
  BUFFD2 U2261 ( .I(completionWriteData_i[0]), .Z(n3141) );
  BUFFD2 U2349 ( .I(completionWriteData_i[55]), .Z(n3196) );
  BUFFD2 U2409 ( .I(completionWriteData_i[61]), .Z(n3202) );
  BUFFD2 U2312 ( .I(completionWriteData_i[36]), .Z(n3177) );
  BUFFD2 U2411 ( .I(completionWriteData_i[63]), .Z(n3204) );
  BUFFD2 U2331 ( .I(completionWriteData_i[53]), .Z(n3194) );
  BUFFD2 U2433 ( .I(completionWriteData_i[67]), .Z(n3208) );
  BUFFD2 U2454 ( .I(completionWriteData_i[69]), .Z(n3210) );
  BUFFD2 U2330 ( .I(completionWriteData_i[52]), .Z(n3193) );
  BUFFD2 U2266 ( .I(completionWriteData_i[5]), .Z(n3146) );
  BUFFD2 U2410 ( .I(completionWriteData_i[62]), .Z(n3203) );
  AOI22D2 U3637 ( .A1(n3297), .A2(\theRegs/completionDataOut[6][2] ), .B1(
        n3703), .B2(\theRegs/completionDataOut[7][2] ), .ZN(n2315) );
  BUFFD2 U2413 ( .I(completionWriteData_i[65]), .Z(n3206) );
  BUFFD2 U2315 ( .I(completionWriteData_i[38]), .Z(n3179) );
  BUFFD2 U2412 ( .I(completionWriteData_i[64]), .Z(n3205) );
  CKBD1 U2326 ( .I(completionWriteData_i[48]), .Z(n3189) );
  BUFFD2 U2414 ( .I(completionWriteData_i[66]), .Z(n3207) );
  BUFFD2 U2437 ( .I(completionWriteData_i[68]), .Z(n3209) );
  ND4D8 U3140 ( .A1(n3047), .A2(n3046), .A3(n3045), .A4(n3044), .ZN(
        decodeReadData2_o[21]) );
  BUFFD2 U2328 ( .I(completionWriteData_i[50]), .Z(n3191) );
  ND4D8 U3851 ( .A1(n2774), .A2(n2773), .A3(n2772), .A4(n2771), .ZN(
        decodeReadData1_o[21]) );
  BUFFD2 U2329 ( .I(completionWriteData_i[51]), .Z(n3192) );
  BUFFD2 U2278 ( .I(completionWriteData_i[12]), .Z(n3153) );
  ND4D8 U3861 ( .A1(n2782), .A2(n2781), .A3(n2780), .A4(n2779), .ZN(
        decodeReadData1_o[19]) );
  BUFFD2 U2279 ( .I(completionWriteData_i[13]), .Z(n3154) );
  AOI22D2 U3457 ( .A1(n3296), .A2(\theRegs/completionDataOut[6][38] ), .B1(
        n4010), .B2(\theRegs/completionDataOut[7][38] ), .ZN(n2459) );
  ND4D8 U3856 ( .A1(n2778), .A2(n2777), .A3(n2776), .A4(n2775), .ZN(
        decodeReadData1_o[20]) );
  AOI22D2 U3452 ( .A1(n3296), .A2(\theRegs/completionDataOut[6][39] ), .B1(
        n4010), .B2(\theRegs/completionDataOut[7][39] ), .ZN(n2463) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[16].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][16] ) );
  AOI22D2 U3472 ( .A1(n3296), .A2(\theRegs/completionDataOut[6][35] ), .B1(
        n4036), .B2(\theRegs/completionDataOut[7][35] ), .ZN(n2447) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[17].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][17] ) );
  BUFFD2 U2281 ( .I(completionWriteData_i[14]), .Z(n3155) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[13].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][13] ) );
  BUFFD2 U2282 ( .I(completionWriteData_i[15]), .Z(n3156) );
  BUFFD1 U2399 ( .I(completionWriteData_i[58]), .Z(n3199) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[16].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][16] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[15].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][15] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[17].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][17] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[19].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][19] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[14].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][14] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[15].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][15] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[18].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][18] ) );
  BUFFD2 U2304 ( .I(completionWriteData_i[30]), .Z(n3171) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[17].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][17] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[14].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][14] ) );
  BUFFD1 U2400 ( .I(completionWriteData_i[59]), .Z(n3200) );
  BUFFD2 U2284 ( .I(completionWriteData_i[16]), .Z(n3157) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[18].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][18] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[19].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][19] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[19].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][19] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[12].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][12] ) );
  BUFFD2 U2285 ( .I(completionWriteData_i[17]), .Z(n3158) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[18].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][18] ) );
  BUFFD2 U2305 ( .I(completionWriteData_i[31]), .Z(n3172) );
  BUFFD2 U2306 ( .I(completionWriteData_i[32]), .Z(n3173) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[21].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][21] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[18].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][18] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[20].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][20] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[21].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][21] ) );
  BUFFD2 U2307 ( .I(completionWriteData_i[33]), .Z(n3174) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[20].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][20] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[13].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][13] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[19].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][19] ) );
  BUFFD2 U2290 ( .I(completionWriteData_i[19]), .Z(n3160) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[21].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][21] ) );
  BUFFD1 U2560 ( .I(decodeWriteData_i[6]), .Z(n3222) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[11].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][11] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[11].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][11] ) );
  BUFFD1 U2521 ( .I(decodeWriteData_i[4]), .Z(n3220) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[11].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][11] ) );
  BUFFD2 U2598 ( .I(decodeReadAddr1_i[0]), .Z(n3231) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[54].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][54] ) );
  AOI22D2 U3104 ( .A1(n2207), .A2(n3240), .B1(n3283), .B2(n3242), .ZN(n2204)
         );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[56].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][56] ) );
  DFQD2 \headTailManager/head_reg[0]  ( .D(n1406), .CP(clk_i), .Q(head[0]) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[20].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][20] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][0] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[57].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][57] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[54].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][54] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[56].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][56] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[21].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][21] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[10].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][10] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[49].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][49] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][6] ) );
  NR4D8 U4176 ( .A1(n3284), .A2(n2221), .A3(n2220), .A4(n2223), .ZN(n2226) );
  BUFFD6 U3062 ( .I(n2584), .Z(n3301) );
  NR3D2 U4188 ( .A1(n3246), .A2(n3243), .A3(n4030), .ZN(n2586) );
  AOI22D4 U3102 ( .A1(tail[0]), .A2(n3239), .B1(tailReset), .B2(n3238), .ZN(
        n4118) );
  NR4D8 U3003 ( .A1(n3212), .A2(n3214), .A3(n3215), .A4(n3211), .ZN(n2177) );
  INR4D2 U2500 ( .A1(n3215), .B1(n3751), .B2(n3211), .B3(n3213), .ZN(n2186) );
  NR4D8 U2416 ( .A1(n3751), .A2(n3851), .A3(n3211), .A4(n3213), .ZN(n2200) );
  NR3D3 U4190 ( .A1(n3246), .A2(n3244), .A3(n3884), .ZN(n2588) );
  INR4D2 U2868 ( .A1(n3751), .B1(n3851), .B2(n3211), .B3(n3212), .ZN(n2195) );
  NR3D3 U4185 ( .A1(n3244), .A2(n3245), .A3(n4009), .ZN(n2587) );
  AOI22D4 U4832 ( .A1(tailReset), .A2(n3285), .B1(n2265), .B2(n3239), .ZN(
        n2227) );
  AO21D4 U2280 ( .A1(n3140), .A2(n3291), .B(reset_i), .Z(n2236) );
  NR3D2 U4153 ( .A1(n3229), .A2(n3225), .A3(n3228), .ZN(n3130) );
  INR4D2 U2667 ( .A1(n3214), .B1(n3851), .B2(n3211), .B3(n3213), .ZN(n2192) );
  NR3D4 U4183 ( .A1(n3243), .A2(n3245), .A3(n4030), .ZN(n2585) );
  IOA21D2 U3014 ( .A1(n3140), .A2(head_o[3]), .B(n2260), .ZN(n2209) );
  INR4D2 U2919 ( .A1(n3851), .B1(n3751), .B2(n3211), .B3(n3212), .ZN(n2189) );
  AOI22D2 U3254 ( .A1(\theRegs/managementDataOut[1][8] ), .A2(n3291), .B1(
        n3276), .B2(\theRegs/managementDataOut[0][8] ), .ZN(n2305) );
  AOI22D2 U3184 ( .A1(\theRegs/completionDataOut[2][13] ), .A2(n3251), .B1(
        \theRegs/completionDataOut[0][13] ), .B2(n3259), .ZN(n3079) );
  AOI22D2 U3239 ( .A1(\theRegs/completionDataOut[2][2] ), .A2(n3252), .B1(
        \theRegs/completionDataOut[0][2] ), .B2(n3260), .ZN(n3123) );
  AOI22D2 U4015 ( .A1(\theRegs/completionDataOut[2][43] ), .A2(n3252), .B1(
        \theRegs/completionDataOut[0][43] ), .B2(n3260), .ZN(n2959) );
  AOI22D2 U3194 ( .A1(\theRegs/completionDataOut[2][11] ), .A2(n3251), .B1(
        \theRegs/completionDataOut[0][11] ), .B2(n3259), .ZN(n3087) );
  AOI22D2 U3229 ( .A1(\theRegs/completionDataOut[2][4] ), .A2(n3252), .B1(
        \theRegs/completionDataOut[0][4] ), .B2(n3260), .ZN(n3115) );
  AOI22D2 U3204 ( .A1(\theRegs/completionDataOut[2][9] ), .A2(n3252), .B1(
        \theRegs/completionDataOut[0][9] ), .B2(n3260), .ZN(n3095) );
  AOI22D2 U3244 ( .A1(\theRegs/completionDataOut[2][1] ), .A2(n3578), .B1(
        \theRegs/completionDataOut[0][1] ), .B2(n3538), .ZN(n3127) );
  AOI22D2 U3224 ( .A1(\theRegs/completionDataOut[2][5] ), .A2(n3578), .B1(
        \theRegs/completionDataOut[0][5] ), .B2(n3538), .ZN(n3111) );
  AOI22D2 U4113 ( .A1(\theRegs/completionDataOut[5][2] ), .A2(n3265), .B1(
        \theRegs/completionDataOut[4][2] ), .B2(n3257), .ZN(n2848) );
  BUFFD1 U2571 ( .I(decodeWriteData_i[8]), .Z(n3224) );
  BUFFD2 U2534 ( .I(decodeWriteData_i[5]), .Z(n3221) );
  AOI22D2 U3853 ( .A1(\theRegs/completionDataOut[5][21] ), .A2(n3265), .B1(
        \theRegs/completionDataOut[4][21] ), .B2(n3257), .ZN(n2772) );
  AOI22D2 U3179 ( .A1(\theRegs/completionDataOut[2][14] ), .A2(n3251), .B1(
        \theRegs/completionDataOut[0][14] ), .B2(n3259), .ZN(n3075) );
  AOI22D2 U3189 ( .A1(\theRegs/completionDataOut[2][12] ), .A2(n3251), .B1(
        \theRegs/completionDataOut[0][12] ), .B2(n3259), .ZN(n3083) );
  AOI22D2 U3214 ( .A1(\theRegs/completionDataOut[2][7] ), .A2(n3578), .B1(
        \theRegs/completionDataOut[0][7] ), .B2(n3538), .ZN(n3103) );
  AOI22D2 U3404 ( .A1(n3294), .A2(\theRegs/completionDataOut[2][49] ), .B1(
        n3289), .B2(\theRegs/completionDataOut[1][49] ), .ZN(n2505) );
  AOI22D2 U4020 ( .A1(\theRegs/completionDataOut[2][44] ), .A2(n3684), .B1(
        \theRegs/completionDataOut[0][44] ), .B2(n3639), .ZN(n2955) );
  AOI22D2 U3169 ( .A1(\theRegs/completionDataOut[2][16] ), .A2(n3251), .B1(
        \theRegs/completionDataOut[0][16] ), .B2(n3259), .ZN(n3067) );
  AOI22D2 U3838 ( .A1(\theRegs/completionDataOut[5][24] ), .A2(n3265), .B1(
        \theRegs/completionDataOut[4][24] ), .B2(n3257), .ZN(n2760) );
  AOI22D2 U3858 ( .A1(\theRegs/completionDataOut[5][20] ), .A2(n3265), .B1(
        \theRegs/completionDataOut[4][20] ), .B2(n3440), .ZN(n2776) );
  AOI22D2 U4090 ( .A1(\theRegs/completionDataOut[2][42] ), .A2(n3684), .B1(
        \theRegs/completionDataOut[0][42] ), .B2(n3639), .ZN(n2963) );
  AOI22D2 U3938 ( .A1(\theRegs/completionDataOut[5][4] ), .A2(n3414), .B1(
        \theRegs/completionDataOut[4][4] ), .B2(n3440), .ZN(n2840) );
  BUFFD1 U2495 ( .I(decodeWriteData_i[0]), .Z(n3216) );
  AOI22D2 U3209 ( .A1(\theRegs/completionDataOut[2][8] ), .A2(n3684), .B1(
        \theRegs/completionDataOut[0][8] ), .B2(n3639), .ZN(n3099) );
  AOI22D2 U3708 ( .A1(\theRegs/completionDataOut[5][51] ), .A2(n3266), .B1(
        \theRegs/completionDataOut[4][51] ), .B2(n3258), .ZN(n2652) );
  AOI22D2 U3913 ( .A1(\theRegs/completionDataOut[5][9] ), .A2(n3414), .B1(
        \theRegs/completionDataOut[4][9] ), .B2(n3440), .ZN(n2820) );
  AOI22D2 U3993 ( .A1(\theRegs/completionDataOut[6][39] ), .A2(n3254), .B1(
        \theRegs/completionDataOut[5][39] ), .B2(n3256), .ZN(n2973) );
  AOI22D2 U4108 ( .A1(\theRegs/completionDataOut[5][1] ), .A2(n3414), .B1(
        \theRegs/completionDataOut[4][1] ), .B2(n3524), .ZN(n2852) );
  AOI22D2 U3199 ( .A1(\theRegs/completionDataOut[2][10] ), .A2(n3684), .B1(
        \theRegs/completionDataOut[0][10] ), .B2(n3639), .ZN(n3091) );
  AOI22D2 U4055 ( .A1(\theRegs/completionDataOut[2][51] ), .A2(n3503), .B1(
        \theRegs/completionDataOut[0][51] ), .B2(n3442), .ZN(n2927) );
  AOI22D2 U3219 ( .A1(\theRegs/completionDataOut[2][6] ), .A2(n3684), .B1(
        \theRegs/completionDataOut[0][6] ), .B2(n3639), .ZN(n3107) );
  AOI22D2 U3893 ( .A1(\theRegs/completionDataOut[5][13] ), .A2(n3414), .B1(
        \theRegs/completionDataOut[4][13] ), .B2(n3524), .ZN(n2804) );
  AOI22D2 U4138 ( .A1(\theRegs/completionDataOut[2][63] ), .A2(n3708), .B1(
        \theRegs/completionDataOut[0][63] ), .B2(n3660), .ZN(n2879) );
  AOI22D2 U3429 ( .A1(n3294), .A2(\theRegs/completionDataOut[2][44] ), .B1(
        n3290), .B2(\theRegs/completionDataOut[1][44] ), .ZN(n2485) );
  AOI22D2 U3908 ( .A1(\theRegs/completionDataOut[5][10] ), .A2(n3434), .B1(
        \theRegs/completionDataOut[4][10] ), .B2(n3524), .ZN(n2816) );
  AOI22D2 U3234 ( .A1(\theRegs/completionDataOut[2][3] ), .A2(n3708), .B1(
        \theRegs/completionDataOut[0][3] ), .B2(n3660), .ZN(n3119) );
  AOI22D2 U3484 ( .A1(n3293), .A2(\theRegs/completionDataOut[2][33] ), .B1(
        n3289), .B2(\theRegs/completionDataOut[1][33] ), .ZN(n2441) );
  AOI22D2 U3933 ( .A1(\theRegs/completionDataOut[5][5] ), .A2(n3434), .B1(
        \theRegs/completionDataOut[4][5] ), .B2(n3524), .ZN(n2836) );
  AOI22D2 U3833 ( .A1(\theRegs/completionDataOut[5][25] ), .A2(n3434), .B1(
        \theRegs/completionDataOut[4][25] ), .B2(n3524), .ZN(n2756) );
  BUFFD1 U2497 ( .I(decodeWriteData_i[2]), .Z(n3218) );
  AOI22D2 U3978 ( .A1(\theRegs/completionDataOut[6][37] ), .A2(n3254), .B1(
        \theRegs/completionDataOut[5][37] ), .B2(n3256), .ZN(n2981) );
  AOI22D2 U3973 ( .A1(\theRegs/completionDataOut[6][36] ), .A2(n3254), .B1(
        \theRegs/completionDataOut[5][36] ), .B2(n3256), .ZN(n2985) );
  AOI22D2 U3998 ( .A1(\theRegs/completionDataOut[6][40] ), .A2(n3254), .B1(
        \theRegs/completionDataOut[5][40] ), .B2(n3256), .ZN(n2969) );
  AOI22D2 U3409 ( .A1(n3850), .A2(\theRegs/completionDataOut[2][48] ), .B1(
        n3290), .B2(\theRegs/completionDataOut[1][48] ), .ZN(n2501) );
  AOI22D2 U3424 ( .A1(n3850), .A2(\theRegs/completionDataOut[2][45] ), .B1(
        n3290), .B2(\theRegs/completionDataOut[1][45] ), .ZN(n2489) );
  AOI22D2 U3247 ( .A1(\theRegs/completionDataOut[6][0] ), .A2(n3253), .B1(
        \theRegs/completionDataOut[5][0] ), .B2(n3255), .ZN(n3137) );
  AOI22D2 U3923 ( .A1(\theRegs/completionDataOut[5][7] ), .A2(n3434), .B1(
        \theRegs/completionDataOut[4][7] ), .B2(n3533), .ZN(n2828) );
  AOI22D2 U4060 ( .A1(\theRegs/completionDataOut[2][52] ), .A2(n3503), .B1(
        \theRegs/completionDataOut[0][52] ), .B2(n3442), .ZN(n2923) );
  AOI22D2 U3988 ( .A1(\theRegs/completionDataOut[6][38] ), .A2(n3254), .B1(
        \theRegs/completionDataOut[5][38] ), .B2(n3256), .ZN(n2977) );
  AOI22D2 U3174 ( .A1(\theRegs/completionDataOut[2][15] ), .A2(n3503), .B1(
        \theRegs/completionDataOut[0][15] ), .B2(n3442), .ZN(n3071) );
  AOI22D2 U3127 ( .A1(\theRegs/completionDataOut[6][24] ), .A2(n3253), .B1(
        \theRegs/completionDataOut[5][24] ), .B2(n3255), .ZN(n3033) );
  AOI22D2 U3888 ( .A1(\theRegs/completionDataOut[5][14] ), .A2(n3486), .B1(
        \theRegs/completionDataOut[4][14] ), .B2(n3533), .ZN(n2800) );
  AOI22D2 U3137 ( .A1(\theRegs/completionDataOut[6][22] ), .A2(n3253), .B1(
        \theRegs/completionDataOut[5][22] ), .B2(n3255), .ZN(n3041) );
  AOI22D2 U3928 ( .A1(\theRegs/completionDataOut[5][6] ), .A2(n3486), .B1(
        \theRegs/completionDataOut[4][6] ), .B2(n3533), .ZN(n2832) );
  AOI22D2 U3828 ( .A1(\theRegs/completionDataOut[5][26] ), .A2(n3496), .B1(
        \theRegs/completionDataOut[4][26] ), .B2(n3533), .ZN(n2752) );
  AOI22D2 U3878 ( .A1(\theRegs/completionDataOut[5][16] ), .A2(n3496), .B1(
        \theRegs/completionDataOut[4][16] ), .B2(n3636), .ZN(n2792) );
  AOI22D2 U3249 ( .A1(\theRegs/completionDataOut[2][0] ), .A2(n3708), .B1(
        \theRegs/completionDataOut[0][0] ), .B2(n3660), .ZN(n3139) );
  AOI22D2 U3883 ( .A1(\theRegs/completionDataOut[5][15] ), .A2(n3496), .B1(
        \theRegs/completionDataOut[4][15] ), .B2(n3636), .ZN(n2796) );
  AOI22D2 U3117 ( .A1(\theRegs/completionDataOut[6][26] ), .A2(n3253), .B1(
        \theRegs/completionDataOut[5][26] ), .B2(n3443), .ZN(n3025) );
  AOI22D2 U3843 ( .A1(\theRegs/completionDataOut[5][23] ), .A2(n3496), .B1(
        \theRegs/completionDataOut[4][23] ), .B2(n3659), .ZN(n2764) );
  AOI22D2 U3713 ( .A1(\theRegs/completionDataOut[5][52] ), .A2(n3266), .B1(
        \theRegs/completionDataOut[4][52] ), .B2(n3258), .ZN(n2648) );
  AOI22D2 U3479 ( .A1(n3292), .A2(\theRegs/completionDataOut[2][34] ), .B1(
        n3290), .B2(\theRegs/completionDataOut[1][34] ), .ZN(n2445) );
  AOI22D2 U3147 ( .A1(\theRegs/completionDataOut[6][20] ), .A2(n3253), .B1(
        \theRegs/completionDataOut[5][20] ), .B2(n3443), .ZN(n3049) );
  AOI22D2 U3142 ( .A1(\theRegs/completionDataOut[6][21] ), .A2(n3476), .B1(
        \theRegs/completionDataOut[5][21] ), .B2(n3443), .ZN(n3045) );
  AOI22D2 U3439 ( .A1(n3850), .A2(\theRegs/completionDataOut[2][42] ), .B1(
        n3290), .B2(\theRegs/completionDataOut[1][42] ), .ZN(n2477) );
  AOI22D2 U3414 ( .A1(n3850), .A2(\theRegs/completionDataOut[2][47] ), .B1(
        n3355), .B2(\theRegs/completionDataOut[1][47] ), .ZN(n2497) );
  AOI22D2 U3863 ( .A1(\theRegs/completionDataOut[5][19] ), .A2(n3496), .B1(
        \theRegs/completionDataOut[4][19] ), .B2(n3659), .ZN(n2780) );
  AOI22D2 U3644 ( .A1(n3292), .A2(\theRegs/completionDataOut[2][1] ), .B1(
        n3291), .B2(\theRegs/completionDataOut[1][1] ), .ZN(n2313) );
  AOI22D2 U3132 ( .A1(\theRegs/completionDataOut[6][23] ), .A2(n3476), .B1(
        \theRegs/completionDataOut[5][23] ), .B2(n3443), .ZN(n3037) );
  AOI22D2 U3474 ( .A1(n3292), .A2(\theRegs/completionDataOut[2][35] ), .B1(
        n3472), .B2(\theRegs/completionDataOut[1][35] ), .ZN(n2449) );
  AOI22D2 U4065 ( .A1(\theRegs/completionDataOut[2][53] ), .A2(n3503), .B1(
        \theRegs/completionDataOut[0][53] ), .B2(n3442), .ZN(n2919) );
  AOI22D2 U3122 ( .A1(\theRegs/completionDataOut[6][25] ), .A2(n3476), .B1(
        \theRegs/completionDataOut[5][25] ), .B2(n3604), .ZN(n3029) );
  AOI22D2 U3970 ( .A1(\theRegs/completionDataOut[2][35] ), .A2(n3708), .B1(
        \theRegs/completionDataOut[0][35] ), .B2(n3660), .ZN(n2991) );
  AOI22D2 U3823 ( .A1(\theRegs/completionDataOut[5][27] ), .A2(n3593), .B1(
        \theRegs/completionDataOut[4][27] ), .B2(n3659), .ZN(n2748) );
  AOI22D2 U4133 ( .A1(\theRegs/completionDataOut[2][62] ), .A2(n3708), .B1(
        \theRegs/completionDataOut[0][62] ), .B2(n3660), .ZN(n2883) );
  AOI22D2 U3703 ( .A1(\theRegs/completionDataOut[5][50] ), .A2(n3266), .B1(
        \theRegs/completionDataOut[4][50] ), .B2(n3258), .ZN(n2656) );
  AOI22D2 U3718 ( .A1(\theRegs/completionDataOut[5][53] ), .A2(n3266), .B1(
        \theRegs/completionDataOut[4][53] ), .B2(n3258), .ZN(n2644) );
  AOI22D2 U3358 ( .A1(\theRegs/completionDataOut[6][28] ), .A2(n3476), .B1(
        \theRegs/completionDataOut[5][28] ), .B2(n3604), .ZN(n3017) );
  AOI22D2 U3202 ( .A1(\theRegs/completionDataOut[6][9] ), .A2(n3522), .B1(
        \theRegs/completionDataOut[5][9] ), .B2(n3604), .ZN(n3093) );
  AOI22D2 U3349 ( .A1(n3926), .A2(\theRegs/completionDataOut[2][59] ), .B1(
        n3355), .B2(\theRegs/completionDataOut[1][59] ), .ZN(n2545) );
  AOI22D2 U3434 ( .A1(n3926), .A2(\theRegs/completionDataOut[2][43] ), .B1(
        n3355), .B2(\theRegs/completionDataOut[1][43] ), .ZN(n2481) );
  BUFFD2 U2496 ( .I(decodeWriteData_i[1]), .Z(n3217) );
  AOI22D2 U3154 ( .A1(\theRegs/completionDataOut[2][19] ), .A2(n3603), .B1(
        \theRegs/completionDataOut[0][19] ), .B2(n3489), .ZN(n3055) );
  AOI22D2 U3918 ( .A1(\theRegs/completionDataOut[5][8] ), .A2(n3617), .B1(
        \theRegs/completionDataOut[4][8] ), .B2(n3659), .ZN(n2824) );
  AOI22D2 U4070 ( .A1(\theRegs/completionDataOut[2][54] ), .A2(n3603), .B1(
        \theRegs/completionDataOut[0][54] ), .B2(n3489), .ZN(n2915) );
  AOI22D2 U4146 ( .A1(\theRegs/completionDataOut[6][61] ), .A2(n3564), .B1(
        \theRegs/completionDataOut[5][61] ), .B2(n3527), .ZN(n2885) );
  AOI22D2 U3898 ( .A1(\theRegs/completionDataOut[5][12] ), .A2(n3617), .B1(
        \theRegs/completionDataOut[4][12] ), .B2(n3773), .ZN(n2808) );
  AOI22D2 U3950 ( .A1(\theRegs/completionDataOut[2][31] ), .A2(n3603), .B1(
        \theRegs/completionDataOut[0][31] ), .B2(n3489), .ZN(n3007) );
  AOI22D2 U3354 ( .A1(n3926), .A2(\theRegs/completionDataOut[2][58] ), .B1(
        n3355), .B2(\theRegs/completionDataOut[1][58] ), .ZN(n2541) );
  AOI22D2 U4085 ( .A1(\theRegs/completionDataOut[2][57] ), .A2(n3621), .B1(
        \theRegs/completionDataOut[0][57] ), .B2(n3507), .ZN(n2903) );
  AOI22D2 U4075 ( .A1(\theRegs/completionDataOut[2][55] ), .A2(n3621), .B1(
        \theRegs/completionDataOut[0][55] ), .B2(n3507), .ZN(n2911) );
  AOI22D2 U3549 ( .A1(n3293), .A2(\theRegs/completionDataOut[2][20] ), .B1(
        n3289), .B2(\theRegs/completionDataOut[1][20] ), .ZN(n2389) );
  AOI22D2 U3149 ( .A1(\theRegs/completionDataOut[2][20] ), .A2(n3621), .B1(
        \theRegs/completionDataOut[0][20] ), .B2(n3507), .ZN(n3051) );
  AOI22D2 U3489 ( .A1(n3293), .A2(\theRegs/completionDataOut[2][32] ), .B1(
        n3289), .B2(\theRegs/completionDataOut[1][32] ), .ZN(n2437) );
  AOI22D2 U4033 ( .A1(\theRegs/completionDataOut[6][47] ), .A2(n3564), .B1(
        \theRegs/completionDataOut[5][47] ), .B2(n3527), .ZN(n2941) );
  AOI22D2 U3242 ( .A1(\theRegs/completionDataOut[6][1] ), .A2(n3522), .B1(
        \theRegs/completionDataOut[5][1] ), .B2(n3604), .ZN(n3125) );
  AOI22D2 U3658 ( .A1(\theRegs/completionDataOut[5][47] ), .A2(n3266), .B1(
        \theRegs/completionDataOut[4][47] ), .B2(n3258), .ZN(n2668) );
  AOI22D2 U4050 ( .A1(\theRegs/completionDataOut[2][50] ), .A2(n3621), .B1(
        \theRegs/completionDataOut[0][50] ), .B2(n3507), .ZN(n2931) );
  AOI22D2 U4040 ( .A1(\theRegs/completionDataOut[2][48] ), .A2(n3621), .B1(
        \theRegs/completionDataOut[0][48] ), .B2(n3507), .ZN(n2939) );
  AOI22D2 U3364 ( .A1(n3926), .A2(\theRegs/completionDataOut[2][57] ), .B1(
        n3355), .B2(\theRegs/completionDataOut[1][57] ), .ZN(n2537) );
  AOI22D2 U3808 ( .A1(\theRegs/completionDataOut[5][30] ), .A2(n3617), .B1(
        \theRegs/completionDataOut[4][30] ), .B2(n3773), .ZN(n2736) );
  AOI22D2 U4118 ( .A1(\theRegs/completionDataOut[5][3] ), .A2(n3617), .B1(
        \theRegs/completionDataOut[4][3] ), .B2(n3773), .ZN(n2844) );
  AOI22D2 U4123 ( .A1(\theRegs/completionDataOut[5][60] ), .A2(n3605), .B1(
        \theRegs/completionDataOut[4][60] ), .B2(n3565), .ZN(n2616) );
  AOI22D2 U3945 ( .A1(\theRegs/completionDataOut[2][30] ), .A2(n3723), .B1(
        \theRegs/completionDataOut[0][30] ), .B2(n3551), .ZN(n3011) );
  AOI22D2 U3768 ( .A1(\theRegs/completionDataOut[5][38] ), .A2(n3605), .B1(
        \theRegs/completionDataOut[4][38] ), .B2(n3565), .ZN(n2704) );
  AO21D4 U2275 ( .A1(n3874), .A2(n3276), .B(reset_i), .Z(n2241) );
  AOI22D2 U4095 ( .A1(\theRegs/completionDataOut[2][58] ), .A2(n3823), .B1(
        \theRegs/completionDataOut[0][58] ), .B2(n3779), .ZN(n2899) );
  AOI22D2 U3965 ( .A1(\theRegs/completionDataOut[2][34] ), .A2(n3723), .B1(
        \theRegs/completionDataOut[0][34] ), .B2(n3551), .ZN(n2995) );
  AOI22D2 U3955 ( .A1(\theRegs/completionDataOut[2][32] ), .A2(n3723), .B1(
        \theRegs/completionDataOut[0][32] ), .B2(n3551), .ZN(n3003) );
  AOI22D2 U3848 ( .A1(\theRegs/completionDataOut[5][22] ), .A2(n3715), .B1(
        \theRegs/completionDataOut[4][22] ), .B2(n3773), .ZN(n2768) );
  AOI22D2 U4038 ( .A1(\theRegs/completionDataOut[6][48] ), .A2(n3564), .B1(
        \theRegs/completionDataOut[5][48] ), .B2(n3527), .ZN(n2937) );
  AOI22D2 U3232 ( .A1(\theRegs/completionDataOut[6][3] ), .A2(n3522), .B1(
        \theRegs/completionDataOut[5][3] ), .B2(n3604), .ZN(n3117) );
  AOI22D2 U4083 ( .A1(\theRegs/completionDataOut[6][57] ), .A2(n3564), .B1(
        \theRegs/completionDataOut[5][57] ), .B2(n3527), .ZN(n2901) );
  AOI22D2 U3953 ( .A1(\theRegs/completionDataOut[6][32] ), .A2(n3522), .B1(
        \theRegs/completionDataOut[5][32] ), .B2(n3616), .ZN(n3001) );
  AOI22D2 U3329 ( .A1(n3926), .A2(\theRegs/completionDataOut[2][63] ), .B1(
        n3371), .B2(\theRegs/completionDataOut[1][63] ), .ZN(n2561) );
  AOI22D2 U4010 ( .A1(\theRegs/completionDataOut[2][29] ), .A2(n3756), .B1(
        \theRegs/completionDataOut[0][29] ), .B2(n3614), .ZN(n3015) );
  AOI22D2 U3968 ( .A1(\theRegs/completionDataOut[6][35] ), .A2(n3564), .B1(
        \theRegs/completionDataOut[5][35] ), .B2(n3527), .ZN(n2989) );
  AOI22D2 U4035 ( .A1(\theRegs/completionDataOut[2][47] ), .A2(n3756), .B1(
        \theRegs/completionDataOut[0][47] ), .B2(n3614), .ZN(n2943) );
  AOI22D2 U3903 ( .A1(\theRegs/completionDataOut[5][11] ), .A2(n3715), .B1(
        \theRegs/completionDataOut[4][11] ), .B2(n3808), .ZN(n2812) );
  AOI22D2 U3399 ( .A1(n3971), .A2(\theRegs/completionDataOut[2][50] ), .B1(
        n3383), .B2(\theRegs/completionDataOut[1][50] ), .ZN(n2509) );
  AOI22D2 U3524 ( .A1(n3293), .A2(\theRegs/completionDataOut[2][25] ), .B1(
        n3289), .B2(\theRegs/completionDataOut[1][25] ), .ZN(n2409) );
  AOI22D2 U4025 ( .A1(\theRegs/completionDataOut[2][45] ), .A2(n3823), .B1(
        \theRegs/completionDataOut[0][45] ), .B2(n3779), .ZN(n2951) );
  AOI22D2 U3773 ( .A1(\theRegs/completionDataOut[5][37] ), .A2(n3605), .B1(
        \theRegs/completionDataOut[4][37] ), .B2(n3565), .ZN(n2708) );
  AOI22D2 U4005 ( .A1(\theRegs/completionDataOut[2][41] ), .A2(n3823), .B1(
        \theRegs/completionDataOut[0][41] ), .B2(n3779), .ZN(n2967) );
  AOI22D2 U4018 ( .A1(\theRegs/completionDataOut[6][44] ), .A2(n3576), .B1(
        \theRegs/completionDataOut[5][44] ), .B2(n3537), .ZN(n2953) );
  AOI22D2 U4141 ( .A1(\theRegs/completionDataOut[6][60] ), .A2(n3576), .B1(
        \theRegs/completionDataOut[5][60] ), .B2(n3537), .ZN(n2889) );
  AOI22D2 U4030 ( .A1(\theRegs/completionDataOut[2][46] ), .A2(n3857), .B1(
        \theRegs/completionDataOut[0][46] ), .B2(n3810), .ZN(n2947) );
  AOI22D2 U4098 ( .A1(\theRegs/completionDataOut[6][64] ), .A2(n3576), .B1(
        \theRegs/completionDataOut[5][64] ), .B2(n3537), .ZN(n2873) );
  AOI22D2 U3980 ( .A1(\theRegs/completionDataOut[2][37] ), .A2(n3857), .B1(
        \theRegs/completionDataOut[0][37] ), .B2(n3810), .ZN(n2983) );
  AOI22D2 U3112 ( .A1(\theRegs/completionDataOut[6][27] ), .A2(n3522), .B1(
        \theRegs/completionDataOut[5][27] ), .B2(n3616), .ZN(n3021) );
  AOI22D2 U3663 ( .A1(\theRegs/completionDataOut[5][46] ), .A2(n3605), .B1(
        \theRegs/completionDataOut[4][46] ), .B2(n3565), .ZN(n2672) );
  AOI22D2 U4063 ( .A1(\theRegs/completionDataOut[6][53] ), .A2(n3576), .B1(
        \theRegs/completionDataOut[5][53] ), .B2(n3537), .ZN(n2917) );
  AOI22D2 U3788 ( .A1(\theRegs/completionDataOut[5][34] ), .A2(n3715), .B1(
        \theRegs/completionDataOut[4][34] ), .B2(n3808), .ZN(n2720) );
  AOI22D2 U4045 ( .A1(\theRegs/completionDataOut[2][49] ), .A2(n3756), .B1(
        \theRegs/completionDataOut[0][49] ), .B2(n3614), .ZN(n2935) );
  AOI22D2 U3960 ( .A1(\theRegs/completionDataOut[2][33] ), .A2(n3756), .B1(
        \theRegs/completionDataOut[0][33] ), .B2(n3614), .ZN(n2999) );
  AOI22D2 U3793 ( .A1(\theRegs/completionDataOut[5][33] ), .A2(n3715), .B1(
        \theRegs/completionDataOut[4][33] ), .B2(n3808), .ZN(n2724) );
  AOI22D2 U3813 ( .A1(\theRegs/completionDataOut[5][29] ), .A2(n3747), .B1(
        \theRegs/completionDataOut[4][29] ), .B2(n3808), .ZN(n2740) );
  AOI22D2 U4080 ( .A1(\theRegs/completionDataOut[2][56] ), .A2(n3863), .B1(
        \theRegs/completionDataOut[0][56] ), .B2(n3669), .ZN(n2907) );
  AOI22D2 U3668 ( .A1(\theRegs/completionDataOut[5][45] ), .A2(n3605), .B1(
        \theRegs/completionDataOut[4][45] ), .B2(n3565), .ZN(n2676) );
  AOI22D2 U4013 ( .A1(\theRegs/completionDataOut[6][43] ), .A2(n3680), .B1(
        \theRegs/completionDataOut[5][43] ), .B2(n3637), .ZN(n2957) );
  AOI22D2 U3162 ( .A1(\theRegs/completionDataOut[6][17] ), .A2(n3552), .B1(
        \theRegs/completionDataOut[5][17] ), .B2(n3616), .ZN(n3061) );
  AOI22D2 U3803 ( .A1(\theRegs/completionDataOut[5][31] ), .A2(n3747), .B1(
        \theRegs/completionDataOut[4][31] ), .B2(n3808), .ZN(n2732) );
  AOI22D2 U3197 ( .A1(\theRegs/completionDataOut[6][10] ), .A2(n3552), .B1(
        \theRegs/completionDataOut[5][10] ), .B2(n3616), .ZN(n3089) );
  AOI22D2 U3778 ( .A1(\theRegs/completionDataOut[5][36] ), .A2(n3611), .B1(
        \theRegs/completionDataOut[4][36] ), .B2(n3577), .ZN(n2712) );
  AOI22D2 U3187 ( .A1(\theRegs/completionDataOut[6][12] ), .A2(n3552), .B1(
        \theRegs/completionDataOut[5][12] ), .B2(n3678), .ZN(n3081) );
  AOI22D2 U3868 ( .A1(\theRegs/completionDataOut[5][18] ), .A2(n3747), .B1(
        \theRegs/completionDataOut[4][18] ), .B2(n3876), .ZN(n2784) );
  AOI22D2 U4143 ( .A1(\theRegs/completionDataOut[2][60] ), .A2(n3857), .B1(
        \theRegs/completionDataOut[0][60] ), .B2(n3810), .ZN(n2891) );
  AOI22D2 U3237 ( .A1(\theRegs/completionDataOut[6][2] ), .A2(n3552), .B1(
        \theRegs/completionDataOut[5][2] ), .B2(n3678), .ZN(n3121) );
  AOI22D2 U3157 ( .A1(\theRegs/completionDataOut[6][18] ), .A2(n3552), .B1(
        \theRegs/completionDataOut[5][18] ), .B2(n3678), .ZN(n3057) );
  AOI22D2 U3738 ( .A1(\theRegs/completionDataOut[5][57] ), .A2(n3611), .B1(
        \theRegs/completionDataOut[4][57] ), .B2(n3577), .ZN(n2628) );
  AOI22D2 U3943 ( .A1(\theRegs/completionDataOut[6][30] ), .A2(n3573), .B1(
        \theRegs/completionDataOut[5][30] ), .B2(n3678), .ZN(n3009) );
  AOI22D2 U3207 ( .A1(\theRegs/completionDataOut[6][8] ), .A2(n3573), .B1(
        \theRegs/completionDataOut[5][8] ), .B2(n3704), .ZN(n3097) );
  AOI22D2 U3212 ( .A1(\theRegs/completionDataOut[6][7] ), .A2(n3573), .B1(
        \theRegs/completionDataOut[5][7] ), .B2(n3704), .ZN(n3101) );
  AOI22D2 U3584 ( .A1(n3293), .A2(\theRegs/completionDataOut[2][13] ), .B1(
        n3664), .B2(\theRegs/completionDataOut[1][13] ), .ZN(n2361) );
  AOI22D2 U4154 ( .A1(\theRegs/completionDataOut[2][59] ), .A2(n3857), .B1(
        \theRegs/completionDataOut[0][59] ), .B2(n3810), .ZN(n2895) );
  AOI22D2 U3419 ( .A1(n3971), .A2(\theRegs/completionDataOut[2][46] ), .B1(
        n3383), .B2(\theRegs/completionDataOut[1][46] ), .ZN(n2493) );
  AOI22D2 U3124 ( .A1(\theRegs/completionDataOut[2][25] ), .A2(n3863), .B1(
        \theRegs/completionDataOut[0][25] ), .B2(n3669), .ZN(n3031) );
  AOI22D2 U3192 ( .A1(\theRegs/completionDataOut[6][11] ), .A2(n3573), .B1(
        \theRegs/completionDataOut[5][11] ), .B2(n3704), .ZN(n3085) );
  AOI22D2 U3139 ( .A1(\theRegs/completionDataOut[2][22] ), .A2(n3863), .B1(
        \theRegs/completionDataOut[0][22] ), .B2(n3669), .ZN(n3043) );
  AOI22D2 U3594 ( .A1(n3501), .A2(\theRegs/completionDataOut[2][11] ), .B1(
        n3664), .B2(\theRegs/completionDataOut[1][11] ), .ZN(n2353) );
  AOI22D2 U3159 ( .A1(\theRegs/completionDataOut[2][18] ), .A2(n3863), .B1(
        \theRegs/completionDataOut[0][18] ), .B2(n3669), .ZN(n3059) );
  AOI22D2 U4148 ( .A1(\theRegs/completionDataOut[2][61] ), .A2(n3857), .B1(
        \theRegs/completionDataOut[0][61] ), .B2(n3810), .ZN(n2887) );
  AOI22D2 U3683 ( .A1(\theRegs/completionDataOut[5][42] ), .A2(n3611), .B1(
        \theRegs/completionDataOut[4][42] ), .B2(n3577), .ZN(n2688) );
  AOI22D2 U3873 ( .A1(\theRegs/completionDataOut[5][17] ), .A2(n3747), .B1(
        \theRegs/completionDataOut[4][17] ), .B2(n3876), .ZN(n2788) );
  AOI22D2 U3222 ( .A1(\theRegs/completionDataOut[6][5] ), .A2(n3819), .B1(
        \theRegs/completionDataOut[5][5] ), .B2(n3704), .ZN(n3109) );
  AOI22D2 U3758 ( .A1(\theRegs/completionDataOut[5][61] ), .A2(n3611), .B1(
        \theRegs/completionDataOut[4][61] ), .B2(n3577), .ZN(n2612) );
  AOI22D2 U3579 ( .A1(n3501), .A2(\theRegs/completionDataOut[2][14] ), .B1(
        n3664), .B2(\theRegs/completionDataOut[1][14] ), .ZN(n2365) );
  AOI22D2 U3114 ( .A1(\theRegs/completionDataOut[2][27] ), .A2(n3891), .B1(
        \theRegs/completionDataOut[0][27] ), .B2(n3738), .ZN(n3023) );
  AOI22D2 U3509 ( .A1(n3501), .A2(\theRegs/completionDataOut[2][28] ), .B1(
        n3664), .B2(\theRegs/completionDataOut[1][28] ), .ZN(n2421) );
  AOI22D2 U3728 ( .A1(\theRegs/completionDataOut[5][55] ), .A2(n3726), .B1(
        \theRegs/completionDataOut[4][55] ), .B2(n3681), .ZN(n2636) );
  AOI22D2 U3182 ( .A1(\theRegs/completionDataOut[6][13] ), .A2(n3819), .B1(
        \theRegs/completionDataOut[5][13] ), .B2(n3704), .ZN(n3077) );
  AOI22D2 U4043 ( .A1(\theRegs/completionDataOut[6][49] ), .A2(n3680), .B1(
        \theRegs/completionDataOut[5][49] ), .B2(n3637), .ZN(n2933) );
  AOI22D2 U3227 ( .A1(\theRegs/completionDataOut[6][4] ), .A2(n3858), .B1(
        \theRegs/completionDataOut[5][4] ), .B2(n3770), .ZN(n3113) );
  AOI22D2 U4088 ( .A1(\theRegs/completionDataOut[6][42] ), .A2(n3680), .B1(
        \theRegs/completionDataOut[5][42] ), .B2(n3637), .ZN(n2961) );
  AOI22D2 U3748 ( .A1(\theRegs/completionDataOut[5][59] ), .A2(n3726), .B1(
        \theRegs/completionDataOut[4][59] ), .B2(n3681), .ZN(n2620) );
  AOI22D2 U3360 ( .A1(\theRegs/completionDataOut[2][28] ), .A2(n3891), .B1(
        \theRegs/completionDataOut[0][28] ), .B2(n3738), .ZN(n3019) );
  AOI22D2 U3723 ( .A1(\theRegs/completionDataOut[5][54] ), .A2(n3726), .B1(
        \theRegs/completionDataOut[4][54] ), .B2(n3681), .ZN(n2640) );
  AOI22D2 U3733 ( .A1(\theRegs/completionDataOut[5][56] ), .A2(n3741), .B1(
        \theRegs/completionDataOut[4][56] ), .B2(n3696), .ZN(n2632) );
  AOI22D2 U3604 ( .A1(n3501), .A2(\theRegs/completionDataOut[2][9] ), .B1(
        n3743), .B2(\theRegs/completionDataOut[1][9] ), .ZN(n2345) );
  AOI22D2 U3108 ( .A1(n3613), .A2(\theRegs/completionDataOut[2][0] ), .B1(
        n3472), .B2(\theRegs/completionDataOut[1][0] ), .ZN(n2309) );
  AOI22D2 U4078 ( .A1(\theRegs/completionDataOut[6][56] ), .A2(n3695), .B1(
        \theRegs/completionDataOut[5][56] ), .B2(n3653), .ZN(n2905) );
  AOI22D2 U3167 ( .A1(\theRegs/completionDataOut[6][16] ), .A2(n3858), .B1(
        \theRegs/completionDataOut[5][16] ), .B2(n3770), .ZN(n3065) );
  AOI22D2 U3152 ( .A1(\theRegs/completionDataOut[6][19] ), .A2(n3858), .B1(
        \theRegs/completionDataOut[5][19] ), .B2(n3770), .ZN(n3053) );
  AOI22D2 U3818 ( .A1(\theRegs/completionDataOut[5][28] ), .A2(n3747), .B1(
        \theRegs/completionDataOut[4][28] ), .B2(n3876), .ZN(n2744) );
  AOI22D2 U3653 ( .A1(\theRegs/completionDataOut[5][48] ), .A2(n3741), .B1(
        \theRegs/completionDataOut[4][48] ), .B2(n3696), .ZN(n2664) );
  AOI22D2 U3177 ( .A1(\theRegs/completionDataOut[6][14] ), .A2(n3858), .B1(
        \theRegs/completionDataOut[5][14] ), .B2(n3799), .ZN(n3073) );
  AOI22D2 U4068 ( .A1(\theRegs/completionDataOut[6][54] ), .A2(n3695), .B1(
        \theRegs/completionDataOut[5][54] ), .B2(n3653), .ZN(n2913) );
  AOI22D2 U3763 ( .A1(\theRegs/completionDataOut[5][62] ), .A2(n3741), .B1(
        \theRegs/completionDataOut[4][62] ), .B2(n3696), .ZN(n2608) );
  AOI22D2 U3983 ( .A1(\theRegs/completionDataOut[5][64] ), .A2(n3866), .B1(
        \theRegs/completionDataOut[4][64] ), .B2(n3822), .ZN(n2600) );
  AOI22D2 U3599 ( .A1(n3501), .A2(\theRegs/completionDataOut[2][10] ), .B1(
        n3743), .B2(\theRegs/completionDataOut[1][10] ), .ZN(n2349) );
  AOI22D2 U3129 ( .A1(\theRegs/completionDataOut[2][24] ), .A2(n3973), .B1(
        \theRegs/completionDataOut[0][24] ), .B2(n3836), .ZN(n3035) );
  AOI22D2 U4058 ( .A1(\theRegs/completionDataOut[6][52] ), .A2(n3695), .B1(
        \theRegs/completionDataOut[5][52] ), .B2(n3653), .ZN(n2921) );
  AOI22D2 U3217 ( .A1(\theRegs/completionDataOut[6][6] ), .A2(n3858), .B1(
        \theRegs/completionDataOut[5][6] ), .B2(n3799), .ZN(n3105) );
  AOI22D2 U4151 ( .A1(\theRegs/completionDataOut[6][59] ), .A2(n3695), .B1(
        \theRegs/completionDataOut[5][59] ), .B2(n3653), .ZN(n2893) );
  AOI22D2 U3698 ( .A1(\theRegs/completionDataOut[5][39] ), .A2(n3866), .B1(
        \theRegs/completionDataOut[4][39] ), .B2(n3822), .ZN(n2700) );
  AOI22D2 U3648 ( .A1(\theRegs/completionDataOut[5][63] ), .A2(n3866), .B1(
        \theRegs/completionDataOut[4][63] ), .B2(n3822), .ZN(n2604) );
  AOI22D2 U3449 ( .A1(n3613), .A2(\theRegs/completionDataOut[2][40] ), .B1(
        n3383), .B2(\theRegs/completionDataOut[1][40] ), .ZN(n2469) );
  AOI22D2 U3172 ( .A1(\theRegs/completionDataOut[6][15] ), .A2(n3858), .B1(
        \theRegs/completionDataOut[5][15] ), .B2(n3799), .ZN(n3069) );
  AOI22D2 U3948 ( .A1(\theRegs/completionDataOut[6][31] ), .A2(n3972), .B1(
        \theRegs/completionDataOut[5][31] ), .B2(n3799), .ZN(n3005) );
  AOI22D2 U3589 ( .A1(n3501), .A2(\theRegs/completionDataOut[2][12] ), .B1(
        n3873), .B2(\theRegs/completionDataOut[1][12] ), .ZN(n2357) );
  AOI22D2 U3673 ( .A1(\theRegs/completionDataOut[5][44] ), .A2(n3892), .B1(
        \theRegs/completionDataOut[4][44] ), .B2(n3847), .ZN(n2680) );
  AOI22D2 U3134 ( .A1(\theRegs/completionDataOut[2][23] ), .A2(n3973), .B1(
        \theRegs/completionDataOut[0][23] ), .B2(n3836), .ZN(n3039) );
  AOI22D2 U3693 ( .A1(\theRegs/completionDataOut[5][40] ), .A2(n3892), .B1(
        \theRegs/completionDataOut[4][40] ), .B2(n3847), .ZN(n2696) );
  AOI22D2 U4008 ( .A1(\theRegs/completionDataOut[6][29] ), .A2(n3972), .B1(
        \theRegs/completionDataOut[5][29] ), .B2(n3929), .ZN(n3013) );
  AOI22D2 U4131 ( .A1(\theRegs/completionDataOut[6][62] ), .A2(n3821), .B1(
        \theRegs/completionDataOut[5][62] ), .B2(n3776), .ZN(n2881) );
  AOI22D2 U3783 ( .A1(\theRegs/completionDataOut[5][35] ), .A2(n3892), .B1(
        \theRegs/completionDataOut[4][35] ), .B2(n3847), .ZN(n2716) );
  AOI22D2 U4073 ( .A1(\theRegs/completionDataOut[6][55] ), .A2(n3821), .B1(
        \theRegs/completionDataOut[5][55] ), .B2(n3776), .ZN(n2909) );
  AOI22D2 U3963 ( .A1(\theRegs/completionDataOut[6][34] ), .A2(n3972), .B1(
        \theRegs/completionDataOut[5][34] ), .B2(n3929), .ZN(n2993) );
  AOI22D2 U3958 ( .A1(\theRegs/completionDataOut[6][33] ), .A2(n3972), .B1(
        \theRegs/completionDataOut[5][33] ), .B2(n3929), .ZN(n2997) );
  AOI22D2 U3798 ( .A1(\theRegs/completionDataOut[5][32] ), .A2(n3928), .B1(
        \theRegs/completionDataOut[4][32] ), .B2(n3876), .ZN(n2728) );
  AOI22D2 U4003 ( .A1(\theRegs/completionDataOut[6][41] ), .A2(n3846), .B1(
        \theRegs/completionDataOut[5][41] ), .B2(n3798), .ZN(n2965) );
  AOI22D2 U3990 ( .A1(\theRegs/completionDataOut[2][38] ), .A2(n3857), .B1(
        \theRegs/completionDataOut[0][38] ), .B2(n3810), .ZN(n2979) );
  AOI22D2 U3624 ( .A1(n3562), .A2(\theRegs/completionDataOut[2][5] ), .B1(
        n3472), .B2(\theRegs/completionDataOut[1][5] ), .ZN(n2329) );
  AOI22D2 U3544 ( .A1(n3568), .A2(\theRegs/completionDataOut[2][21] ), .B1(
        n3873), .B2(\theRegs/completionDataOut[1][21] ), .ZN(n2393) );
  AOI22D2 U3569 ( .A1(n3568), .A2(\theRegs/completionDataOut[2][16] ), .B1(
        n3873), .B2(\theRegs/completionDataOut[1][16] ), .ZN(n2373) );
  AOI22D2 U4048 ( .A1(\theRegs/completionDataOut[6][50] ), .A2(n3846), .B1(
        \theRegs/completionDataOut[5][50] ), .B2(n3798), .ZN(n2929) );
  AOI22D2 U3119 ( .A1(\theRegs/completionDataOut[2][26] ), .A2(n3973), .B1(
        \theRegs/completionDataOut[0][26] ), .B2(n3836), .ZN(n3027) );
  AOI22D2 U4000 ( .A1(\theRegs/completionDataOut[2][40] ), .A2(n3961), .B1(
        \theRegs/completionDataOut[0][40] ), .B2(n3912), .ZN(n2971) );
  AOI22D2 U4028 ( .A1(\theRegs/completionDataOut[6][46] ), .A2(n3846), .B1(
        \theRegs/completionDataOut[5][46] ), .B2(n3798), .ZN(n2945) );
  AOI22D2 U3688 ( .A1(\theRegs/completionDataOut[5][41] ), .A2(n3892), .B1(
        \theRegs/completionDataOut[4][41] ), .B2(n3847), .ZN(n2692) );
  AOI22D2 U3144 ( .A1(\theRegs/completionDataOut[2][21] ), .A2(n3973), .B1(
        \theRegs/completionDataOut[0][21] ), .B2(n3836), .ZN(n3047) );
  AOI22D2 U3619 ( .A1(n3568), .A2(\theRegs/completionDataOut[2][6] ), .B1(
        n3472), .B2(\theRegs/completionDataOut[1][6] ), .ZN(n2333) );
  AOI22D2 U3394 ( .A1(n3971), .A2(\theRegs/completionDataOut[2][51] ), .B1(
        n3383), .B2(\theRegs/completionDataOut[1][51] ), .ZN(n2513) );
  AOI22D2 U4136 ( .A1(\theRegs/completionDataOut[6][63] ), .A2(n3846), .B1(
        \theRegs/completionDataOut[5][63] ), .B2(n3798), .ZN(n2877) );
  AOI22D2 U4100 ( .A1(\theRegs/completionDataOut[2][64] ), .A2(n3961), .B1(
        \theRegs/completionDataOut[0][64] ), .B2(n3912), .ZN(n2875) );
  AOI22D2 U4023 ( .A1(\theRegs/completionDataOut[6][45] ), .A2(n3962), .B1(
        \theRegs/completionDataOut[5][45] ), .B2(n3913), .ZN(n2949) );
  AOI22D2 U3444 ( .A1(n3971), .A2(\theRegs/completionDataOut[2][41] ), .B1(
        n3383), .B2(\theRegs/completionDataOut[1][41] ), .ZN(n2473) );
  AOI22D2 U3975 ( .A1(\theRegs/completionDataOut[2][36] ), .A2(n3961), .B1(
        \theRegs/completionDataOut[0][36] ), .B2(n3912), .ZN(n2987) );
  AOI22D2 U3519 ( .A1(n3568), .A2(\theRegs/completionDataOut[2][26] ), .B1(
        n3873), .B2(\theRegs/completionDataOut[1][26] ), .ZN(n2413) );
  AOI22D2 U3164 ( .A1(\theRegs/completionDataOut[2][17] ), .A2(n3973), .B1(
        \theRegs/completionDataOut[0][17] ), .B2(n3836), .ZN(n3063) );
  AOI22D2 U3514 ( .A1(n3634), .A2(\theRegs/completionDataOut[2][27] ), .B1(
        n3927), .B2(\theRegs/completionDataOut[1][27] ), .ZN(n2417) );
  AOI22D2 U3504 ( .A1(n3634), .A2(\theRegs/completionDataOut[2][29] ), .B1(
        n3927), .B2(\theRegs/completionDataOut[1][29] ), .ZN(n2425) );
  AOI22D2 U3678 ( .A1(\theRegs/completionDataOut[5][43] ), .A2(n3892), .B1(
        \theRegs/completionDataOut[4][43] ), .B2(n3847), .ZN(n2684) );
  AOI22D2 U3499 ( .A1(n3647), .A2(\theRegs/completionDataOut[2][30] ), .B1(
        n3927), .B2(\theRegs/completionDataOut[1][30] ), .ZN(n2429) );
  AOI22D2 U3529 ( .A1(n3647), .A2(\theRegs/completionDataOut[2][24] ), .B1(
        n3927), .B2(\theRegs/completionDataOut[1][24] ), .ZN(n2405) );
  AOI22D2 U3344 ( .A1(n3971), .A2(\theRegs/completionDataOut[2][60] ), .B1(
        n3396), .B2(\theRegs/completionDataOut[1][60] ), .ZN(n2549) );
  AOI22D2 U4093 ( .A1(\theRegs/completionDataOut[6][58] ), .A2(n3962), .B1(
        \theRegs/completionDataOut[5][58] ), .B2(n3913), .ZN(n2897) );
  AOI22D2 U3384 ( .A1(n3971), .A2(\theRegs/completionDataOut[2][53] ), .B1(
        n3396), .B2(\theRegs/completionDataOut[1][53] ), .ZN(n2521) );
  AOI22D2 U3753 ( .A1(\theRegs/completionDataOut[5][49] ), .A2(n3992), .B1(
        \theRegs/completionDataOut[4][49] ), .B2(n3963), .ZN(n2660) );
  AOI22D2 U3369 ( .A1(n3993), .A2(\theRegs/completionDataOut[2][56] ), .B1(
        n3396), .B2(\theRegs/completionDataOut[1][56] ), .ZN(n2533) );
  AOI22D2 U3559 ( .A1(n3647), .A2(\theRegs/completionDataOut[2][18] ), .B1(
        n3927), .B2(\theRegs/completionDataOut[1][18] ), .ZN(n2381) );
  AOI22D2 U3334 ( .A1(n3613), .A2(\theRegs/completionDataOut[2][62] ), .B1(
        n3396), .B2(\theRegs/completionDataOut[1][62] ), .ZN(n2557) );
  AOI22D2 U4053 ( .A1(\theRegs/completionDataOut[6][51] ), .A2(n3962), .B1(
        \theRegs/completionDataOut[5][51] ), .B2(n3913), .ZN(n2925) );
  AOI22D2 U3554 ( .A1(n3647), .A2(\theRegs/completionDataOut[2][19] ), .B1(
        n3927), .B2(\theRegs/completionDataOut[1][19] ), .ZN(n2385) );
  AOI22D2 U3574 ( .A1(n3647), .A2(\theRegs/completionDataOut[2][15] ), .B1(
        n3965), .B2(\theRegs/completionDataOut[1][15] ), .ZN(n2369) );
  AOI22D2 U3324 ( .A1(n3731), .A2(\theRegs/completionDataOut[2][64] ), .B1(
        n3396), .B2(\theRegs/completionDataOut[1][64] ), .ZN(n2565) );
  AOI22D2 U3995 ( .A1(\theRegs/completionDataOut[2][39] ), .A2(n3961), .B1(
        \theRegs/completionDataOut[0][39] ), .B2(n3912), .ZN(n2975) );
  AOI22D2 U4103 ( .A1(\theRegs/completionDataOut[5][0] ), .A2(n3928), .B1(
        \theRegs/completionDataOut[4][0] ), .B2(n3876), .ZN(n2864) );
  AOI22D2 U3743 ( .A1(\theRegs/completionDataOut[5][58] ), .A2(n3992), .B1(
        \theRegs/completionDataOut[4][58] ), .B2(n3963), .ZN(n2624) );
  AOI22D2 U3379 ( .A1(n3993), .A2(\theRegs/completionDataOut[2][54] ), .B1(
        n3419), .B2(\theRegs/completionDataOut[1][54] ), .ZN(n2525) );
  AOI22D2 U3494 ( .A1(n3721), .A2(\theRegs/completionDataOut[2][31] ), .B1(
        n3965), .B2(\theRegs/completionDataOut[1][31] ), .ZN(n2433) );
  AOI22D2 U3534 ( .A1(n3737), .A2(\theRegs/completionDataOut[2][23] ), .B1(
        n3965), .B2(\theRegs/completionDataOut[1][23] ), .ZN(n2401) );
  AOI22D2 U3389 ( .A1(n3993), .A2(\theRegs/completionDataOut[2][52] ), .B1(
        n3419), .B2(\theRegs/completionDataOut[1][52] ), .ZN(n2517) );
  AOI22D2 U3609 ( .A1(n3737), .A2(\theRegs/completionDataOut[2][8] ), .B1(
        n3472), .B2(\theRegs/completionDataOut[1][8] ), .ZN(n2341) );
  AOI22D2 U3374 ( .A1(n3993), .A2(\theRegs/completionDataOut[2][55] ), .B1(
        n3419), .B2(\theRegs/completionDataOut[1][55] ), .ZN(n2529) );
  AOI22D2 U3564 ( .A1(n3737), .A2(\theRegs/completionDataOut[2][17] ), .B1(
        n3965), .B2(\theRegs/completionDataOut[1][17] ), .ZN(n2377) );
  AOI22D2 U3339 ( .A1(n3993), .A2(\theRegs/completionDataOut[2][61] ), .B1(
        n3429), .B2(\theRegs/completionDataOut[1][61] ), .ZN(n2553) );
  AOI22D2 U3539 ( .A1(n3737), .A2(\theRegs/completionDataOut[2][22] ), .B1(
        n3965), .B2(\theRegs/completionDataOut[1][22] ), .ZN(n2397) );
  AOI22D2 U3469 ( .A1(n3731), .A2(\theRegs/completionDataOut[2][36] ), .B1(
        n3607), .B2(\theRegs/completionDataOut[1][36] ), .ZN(n2453) );
  AOI22D2 U3629 ( .A1(n3813), .A2(\theRegs/completionDataOut[2][4] ), .B1(
        n3607), .B2(\theRegs/completionDataOut[1][4] ), .ZN(n2325) );
  ND2D1 U3250 ( .A1(n2247), .A2(n4028), .ZN(nextTail_o[1]) );
  AOI22D2 U3464 ( .A1(n3731), .A2(\theRegs/completionDataOut[2][37] ), .B1(
        n3607), .B2(\theRegs/completionDataOut[1][37] ), .ZN(n2457) );
  AOI22D2 U3639 ( .A1(n3731), .A2(\theRegs/completionDataOut[2][2] ), .B1(
        n3607), .B2(\theRegs/completionDataOut[1][2] ), .ZN(n2317) );
  AOI22D2 U3454 ( .A1(n3731), .A2(\theRegs/completionDataOut[2][39] ), .B1(
        n3607), .B2(\theRegs/completionDataOut[1][39] ), .ZN(n2465) );
  AOI22D2 U3298 ( .A1(n3286), .A2(\theRegs/completionDataOut[3][69] ), .B1(
        n3755), .B2(\theRegs/completionDataOut[2][69] ), .ZN(n2591) );
  NR3D1 U4838 ( .A1(n3284), .A2(n3887), .A3(n2220), .ZN(n2224) );
  IND2D2 U4827 ( .A1(n2246), .B1(n2243), .ZN(n2237) );
  OAI22D2 U4157 ( .A1(n4041), .A2(n2257), .B1(n2256), .B2(n3307), .ZN(n1404)
         );
  CKND2 U3103 ( .I(updateTail_i), .ZN(n2269) );
  AOI22D4 U4194 ( .A1(tail[0]), .A2(n2262), .B1(tail[1]), .B2(n3238), .ZN(
        n2263) );
  AOI22D2 U4844 ( .A1(n3247), .A2(n4007), .B1(n2256), .B2(n3250), .ZN(n1406)
         );
  AOI22D4 U4840 ( .A1(n3241), .A2(n3245), .B1(n3246), .B2(n4011), .ZN(
        head_o[1]) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][3] ) );
  BUFFD2 U2563 ( .I(decodeWriteData_i[7]), .Z(n3223) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][0] ) );
  ND2D1 U4169 ( .A1(n2268), .A2(\add_x_6/n1 ), .ZN(n2208) );
  BUFFD2 U2594 ( .I(decodeReadAddr2_i[1]), .Z(n3227) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[38].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][38] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][2] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[39].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][39] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][7] ) );
  NR3D1 U4128 ( .A1(n3233), .A2(n3234), .A3(n3232), .ZN(n3736) );
  NR3D1 U4155 ( .A1(n3229), .A2(n3227), .A3(n3226), .ZN(n3839) );
  AOI22D4 U3101 ( .A1(tailReset), .A2(n3983), .B1(n2262), .B2(n3239), .ZN(
        n2221) );
  AOI221D4 U2287 ( .A1(n3247), .A2(tail[0]), .B1(head_o[0]), .B2(n3238), .C(
        n2206), .ZN(n2270) );
  ND4D8 U3466 ( .A1(n2454), .A2(n2453), .A3(n2452), .A4(n2451), .ZN(
        commitReadData_o[36]) );
  ND4D8 U3461 ( .A1(n2458), .A2(n2457), .A3(n2456), .A4(n2455), .ZN(
        commitReadData_o[37]) );
  AOI31D4 U4181 ( .A1(n2243), .A2(nextTail_o[0]), .A3(n3305), .B(n2241), .ZN(
        n2244) );
  NR2D3 U4823 ( .A1(n2232), .A2(n2233), .ZN(n2235) );
  ND4D8 U3451 ( .A1(n2466), .A2(n2465), .A3(n2464), .A4(n2463), .ZN(
        commitReadData_o[39]) );
  NR3D2 U4200 ( .A1(n3233), .A2(n3232), .A3(n3235), .ZN(n2859) );
  BUFFD2 U2665 ( .I(head[1]), .Z(n3243) );
  ND4D8 U3621 ( .A1(n2330), .A2(n2329), .A3(n2328), .A4(n2327), .ZN(
        commitReadData_o[5]) );
  ND4D8 U3251 ( .A1(n2306), .A2(n2305), .A3(n2304), .A4(n2303), .ZN(
        commitReadData_o[78]) );
  ND4D3 U3301 ( .A1(n2582), .A2(n2581), .A3(n2580), .A4(n2579), .ZN(
        commitReadData_o[68]) );
  ND4D3 U3276 ( .A1(n2286), .A2(n2285), .A3(n3936), .A4(n2283), .ZN(
        commitReadData_o[73]) );
  ND4D3 U3271 ( .A1(n2290), .A2(n2289), .A3(n3937), .A4(n2287), .ZN(
        commitReadData_o[74]) );
  ND4D3 U3256 ( .A1(n2302), .A2(n2301), .A3(n3939), .A4(n2299), .ZN(
        commitReadData_o[77]) );
  ND4D3 U3266 ( .A1(n2294), .A2(n2293), .A3(n3938), .A4(n2291), .ZN(
        commitReadData_o[75]) );
  AOI22D2 U3550 ( .A1(n3299), .A2(\theRegs/completionDataOut[4][20] ), .B1(
        n3276), .B2(\theRegs/completionDataOut[0][20] ), .ZN(n2390) );
  ND4D2 U3281 ( .A1(n2282), .A2(n2281), .A3(n2280), .A4(n2279), .ZN(
        commitReadData_o[72]) );
  AOI22D2 U3837 ( .A1(\theRegs/completionDataOut[7][24] ), .A2(n3273), .B1(
        \theRegs/completionDataOut[6][24] ), .B2(n3267), .ZN(n2759) );
  AOI22D2 U3797 ( .A1(\theRegs/completionDataOut[7][32] ), .A2(n3273), .B1(
        \theRegs/completionDataOut[6][32] ), .B2(n3267), .ZN(n2727) );
  AOI22D2 U3116 ( .A1(\theRegs/completionDataOut[7][26] ), .A2(n3281), .B1(
        \theRegs/completionDataOut[4][26] ), .B2(n3269), .ZN(n3024) );
  AOI22D2 U3684 ( .A1(\theRegs/completionDataOut[3][42] ), .A2(n3272), .B1(
        \theRegs/completionDataOut[1][42] ), .B2(n3237), .ZN(n2689) );
  ND3D2 U4184 ( .A1(n2243), .A2(nextTail_o[0]), .A3(n3305), .ZN(n2240) );
  AOI22D2 U4009 ( .A1(\theRegs/completionDataOut[3][29] ), .A2(n3277), .B1(
        \theRegs/completionDataOut[1][29] ), .B2(n3261), .ZN(n3014) );
  AOI22D2 U3525 ( .A1(n3299), .A2(\theRegs/completionDataOut[4][25] ), .B1(
        n3276), .B2(\theRegs/completionDataOut[0][25] ), .ZN(n2410) );
  AOI22D2 U3126 ( .A1(\theRegs/completionDataOut[7][24] ), .A2(n3281), .B1(
        \theRegs/completionDataOut[4][24] ), .B2(n3269), .ZN(n3032) );
  AOI22D2 U3121 ( .A1(\theRegs/completionDataOut[7][25] ), .A2(n3281), .B1(
        \theRegs/completionDataOut[4][25] ), .B2(n3269), .ZN(n3028) );
  AOI22D2 U4132 ( .A1(\theRegs/completionDataOut[3][62] ), .A2(n3278), .B1(
        \theRegs/completionDataOut[1][62] ), .B2(n3262), .ZN(n2882) );
  ND4D8 U3261 ( .A1(n2298), .A2(n2297), .A3(n2296), .A4(n2295), .ZN(
        commitReadData_o[76]) );
  AOI22D2 U3857 ( .A1(\theRegs/completionDataOut[7][20] ), .A2(n3273), .B1(
        \theRegs/completionDataOut[6][20] ), .B2(n3267), .ZN(n2775) );
  AOI22D2 U3527 ( .A1(n3295), .A2(\theRegs/completionDataOut[6][24] ), .B1(
        n3302), .B2(\theRegs/completionDataOut[7][24] ), .ZN(n2403) );
  AOI22D2 U4089 ( .A1(\theRegs/completionDataOut[3][42] ), .A2(n3278), .B1(
        \theRegs/completionDataOut[1][42] ), .B2(n3262), .ZN(n2962) );
  AOI22D2 U3852 ( .A1(\theRegs/completionDataOut[7][21] ), .A2(n3273), .B1(
        \theRegs/completionDataOut[6][21] ), .B2(n3267), .ZN(n2771) );
  AOI22D2 U3547 ( .A1(n3295), .A2(\theRegs/completionDataOut[6][20] ), .B1(
        n3302), .B2(\theRegs/completionDataOut[7][20] ), .ZN(n2387) );
  AOI22D2 U3545 ( .A1(n3299), .A2(\theRegs/completionDataOut[4][21] ), .B1(
        n3276), .B2(\theRegs/completionDataOut[0][21] ), .ZN(n2394) );
  AOI22D2 U3492 ( .A1(n3295), .A2(\theRegs/completionDataOut[6][31] ), .B1(
        n3302), .B2(\theRegs/completionDataOut[7][31] ), .ZN(n2431) );
  AOI22D2 U3952 ( .A1(\theRegs/completionDataOut[7][32] ), .A2(n3281), .B1(
        \theRegs/completionDataOut[4][32] ), .B2(n3269), .ZN(n3000) );
  AOI22D2 U3669 ( .A1(\theRegs/completionDataOut[3][45] ), .A2(n3272), .B1(
        \theRegs/completionDataOut[1][45] ), .B2(n3237), .ZN(n2677) );
  AOI22D2 U3809 ( .A1(\theRegs/completionDataOut[3][30] ), .A2(n3271), .B1(
        \theRegs/completionDataOut[1][30] ), .B2(n3236), .ZN(n2737) );
  AOI22D2 U4022 ( .A1(\theRegs/completionDataOut[7][45] ), .A2(n3282), .B1(
        \theRegs/completionDataOut[4][45] ), .B2(n3270), .ZN(n2948) );
  AOI22D2 U3530 ( .A1(n3344), .A2(\theRegs/completionDataOut[4][24] ), .B1(
        n3356), .B2(\theRegs/completionDataOut[0][24] ), .ZN(n2406) );
  AOI22D2 U3146 ( .A1(\theRegs/completionDataOut[7][20] ), .A2(n3281), .B1(
        \theRegs/completionDataOut[4][20] ), .B2(n3269), .ZN(n3048) );
  AOI22D2 U3487 ( .A1(n3296), .A2(\theRegs/completionDataOut[6][32] ), .B1(
        n3304), .B2(\theRegs/completionDataOut[7][32] ), .ZN(n2435) );
  AOI22D2 U3679 ( .A1(\theRegs/completionDataOut[3][43] ), .A2(n3272), .B1(
        \theRegs/completionDataOut[1][43] ), .B2(n3237), .ZN(n2685) );
  AOI22D2 U3131 ( .A1(\theRegs/completionDataOut[7][23] ), .A2(n3343), .B1(
        \theRegs/completionDataOut[4][23] ), .B2(n3464), .ZN(n3036) );
  AOI22D2 U3814 ( .A1(\theRegs/completionDataOut[3][29] ), .A2(n3271), .B1(
        \theRegs/completionDataOut[1][29] ), .B2(n3236), .ZN(n2741) );
  ND4D2 U3286 ( .A1(n2278), .A2(n2277), .A3(n3934), .A4(n2275), .ZN(
        commitReadData_o[71]) );
  AOI22D2 U3764 ( .A1(\theRegs/completionDataOut[3][62] ), .A2(n3272), .B1(
        \theRegs/completionDataOut[1][62] ), .B2(n3237), .ZN(n2609) );
  ND4D2 U3291 ( .A1(n2274), .A2(n2273), .A3(n3935), .A4(n2271), .ZN(
        commitReadData_o[70]) );
  AOI22D2 U3874 ( .A1(\theRegs/completionDataOut[3][17] ), .A2(n3409), .B1(
        \theRegs/completionDataOut[1][17] ), .B2(n3394), .ZN(n2789) );
  AOI22D2 U3747 ( .A1(\theRegs/completionDataOut[7][59] ), .A2(n3274), .B1(
        \theRegs/completionDataOut[6][59] ), .B2(n3268), .ZN(n2619) );
  AOI22D2 U3141 ( .A1(\theRegs/completionDataOut[7][21] ), .A2(n3343), .B1(
        \theRegs/completionDataOut[4][21] ), .B2(n3464), .ZN(n3044) );
  AOI22D2 U4137 ( .A1(\theRegs/completionDataOut[3][63] ), .A2(n3278), .B1(
        \theRegs/completionDataOut[1][63] ), .B2(n3262), .ZN(n2878) );
  AOI22D2 U3794 ( .A1(\theRegs/completionDataOut[3][33] ), .A2(n3409), .B1(
        \theRegs/completionDataOut[1][33] ), .B2(n3394), .ZN(n2725) );
  AOI22D2 U3804 ( .A1(\theRegs/completionDataOut[3][31] ), .A2(n3409), .B1(
        \theRegs/completionDataOut[1][31] ), .B2(n3394), .ZN(n2733) );
  AOI22D2 U4147 ( .A1(\theRegs/completionDataOut[3][61] ), .A2(n3278), .B1(
        \theRegs/completionDataOut[1][61] ), .B2(n3262), .ZN(n2886) );
  AOI22D2 U3989 ( .A1(\theRegs/completionDataOut[3][38] ), .A2(n3439), .B1(
        \theRegs/completionDataOut[1][38] ), .B2(n3408), .ZN(n2978) );
  AOI22D2 U3844 ( .A1(\theRegs/completionDataOut[3][23] ), .A2(n3409), .B1(
        \theRegs/completionDataOut[1][23] ), .B2(n3394), .ZN(n2765) );
  AOI22D2 U3849 ( .A1(\theRegs/completionDataOut[3][22] ), .A2(n3437), .B1(
        \theRegs/completionDataOut[1][22] ), .B2(n3406), .ZN(n2769) );
  AOI22D2 U3585 ( .A1(n3344), .A2(\theRegs/completionDataOut[4][13] ), .B1(
        n3356), .B2(\theRegs/completionDataOut[0][13] ), .ZN(n2362) );
  AOI22D2 U3497 ( .A1(n3295), .A2(\theRegs/completionDataOut[6][30] ), .B1(
        n3302), .B2(\theRegs/completionDataOut[7][30] ), .ZN(n2427) );
  AOI22D2 U4142 ( .A1(\theRegs/completionDataOut[3][60] ), .A2(n3439), .B1(
        \theRegs/completionDataOut[1][60] ), .B2(n3408), .ZN(n2890) );
  AOI22D2 U3535 ( .A1(n3344), .A2(\theRegs/completionDataOut[4][23] ), .B1(
        n3356), .B2(\theRegs/completionDataOut[0][23] ), .ZN(n2402) );
  AOI22D2 U4047 ( .A1(\theRegs/completionDataOut[7][50] ), .A2(n3282), .B1(
        \theRegs/completionDataOut[4][50] ), .B2(n3270), .ZN(n2928) );
  AOI22D2 U3532 ( .A1(n3295), .A2(\theRegs/completionDataOut[6][23] ), .B1(
        n3642), .B2(\theRegs/completionDataOut[7][23] ), .ZN(n2399) );
  AOI22D2 U3949 ( .A1(\theRegs/completionDataOut[3][31] ), .A2(n3277), .B1(
        \theRegs/completionDataOut[1][31] ), .B2(n3261), .ZN(n3006) );
  AOI22D2 U3357 ( .A1(\theRegs/completionDataOut[7][28] ), .A2(n3343), .B1(
        \theRegs/completionDataOut[4][28] ), .B2(n3464), .ZN(n3016) );
  AOI22D2 U3542 ( .A1(n3457), .A2(\theRegs/completionDataOut[6][21] ), .B1(
        n3642), .B2(\theRegs/completionDataOut[7][21] ), .ZN(n2391) );
  AOI22D2 U3111 ( .A1(\theRegs/completionDataOut[7][27] ), .A2(n3343), .B1(
        \theRegs/completionDataOut[4][27] ), .B2(n3464), .ZN(n3020) );
  AOI22D2 U3822 ( .A1(\theRegs/completionDataOut[7][27] ), .A2(n3273), .B1(
        \theRegs/completionDataOut[6][27] ), .B2(n3397), .ZN(n2747) );
  AOI22D2 U3799 ( .A1(\theRegs/completionDataOut[3][32] ), .A2(n3437), .B1(
        \theRegs/completionDataOut[1][32] ), .B2(n3406), .ZN(n2729) );
  AOI22D2 U3161 ( .A1(\theRegs/completionDataOut[7][17] ), .A2(n3343), .B1(
        \theRegs/completionDataOut[4][17] ), .B2(n3464), .ZN(n3060) );
  AOI22D2 U3689 ( .A1(\theRegs/completionDataOut[3][41] ), .A2(n3272), .B1(
        \theRegs/completionDataOut[1][41] ), .B2(n3237), .ZN(n2693) );
  AOI22D2 U3133 ( .A1(\theRegs/completionDataOut[3][23] ), .A2(n3277), .B1(
        \theRegs/completionDataOut[1][23] ), .B2(n3261), .ZN(n3038) );
  AOI22D2 U4029 ( .A1(\theRegs/completionDataOut[3][46] ), .A2(n3474), .B1(
        \theRegs/completionDataOut[1][46] ), .B2(n3446), .ZN(n2946) );
  AOI22D2 U3867 ( .A1(\theRegs/completionDataOut[7][18] ), .A2(n3416), .B1(
        \theRegs/completionDataOut[6][18] ), .B2(n3397), .ZN(n2783) );
  AOI22D2 U3156 ( .A1(\theRegs/completionDataOut[7][18] ), .A2(n3346), .B1(
        \theRegs/completionDataOut[4][18] ), .B2(n3523), .ZN(n3056) );
  AOI22D2 U4094 ( .A1(\theRegs/completionDataOut[3][58] ), .A2(n3474), .B1(
        \theRegs/completionDataOut[1][58] ), .B2(n3446), .ZN(n2898) );
  AOI22D2 U3749 ( .A1(\theRegs/completionDataOut[3][59] ), .A2(n3458), .B1(
        \theRegs/completionDataOut[1][59] ), .B2(n3526), .ZN(n2621) );
  AOI22D2 U3802 ( .A1(\theRegs/completionDataOut[7][31] ), .A2(n3416), .B1(
        \theRegs/completionDataOut[6][31] ), .B2(n3397), .ZN(n2731) );
  AOI22D2 U3787 ( .A1(\theRegs/completionDataOut[7][34] ), .A2(n3416), .B1(
        \theRegs/completionDataOut[6][34] ), .B2(n3268), .ZN(n2719) );
  AOI22D2 U3759 ( .A1(\theRegs/completionDataOut[3][61] ), .A2(n3458), .B1(
        \theRegs/completionDataOut[1][61] ), .B2(n3526), .ZN(n2613) );
  AOI22D2 U3842 ( .A1(\theRegs/completionDataOut[7][23] ), .A2(n3416), .B1(
        \theRegs/completionDataOut[6][23] ), .B2(n3397), .ZN(n2763) );
  AOI22D2 U3864 ( .A1(\theRegs/completionDataOut[3][19] ), .A2(n3437), .B1(
        \theRegs/completionDataOut[1][19] ), .B2(n3406), .ZN(n2781) );
  AOI22D2 U3482 ( .A1(n3296), .A2(\theRegs/completionDataOut[6][33] ), .B1(
        n3304), .B2(\theRegs/completionDataOut[7][33] ), .ZN(n2439) );
  AOI22D2 U3734 ( .A1(\theRegs/completionDataOut[3][56] ), .A2(n3458), .B1(
        \theRegs/completionDataOut[1][56] ), .B2(n3526), .ZN(n2633) );
  AOI22D2 U3138 ( .A1(\theRegs/completionDataOut[3][22] ), .A2(n3277), .B1(
        \theRegs/completionDataOut[1][22] ), .B2(n3261), .ZN(n3042) );
  AOI22D2 U3590 ( .A1(n3344), .A2(\theRegs/completionDataOut[4][12] ), .B1(
        n3356), .B2(\theRegs/completionDataOut[0][12] ), .ZN(n2358) );
  AOI22D2 U4049 ( .A1(\theRegs/completionDataOut[3][50] ), .A2(n3474), .B1(
        \theRegs/completionDataOut[1][50] ), .B2(n3446), .ZN(n2930) );
  AOI22D2 U4024 ( .A1(\theRegs/completionDataOut[3][45] ), .A2(n3474), .B1(
        \theRegs/completionDataOut[1][45] ), .B2(n3446), .ZN(n2950) );
  AOI22D2 U3704 ( .A1(\theRegs/completionDataOut[3][50] ), .A2(n3458), .B1(
        \theRegs/completionDataOut[1][50] ), .B2(n3526), .ZN(n2657) );
  AOI22D2 U4004 ( .A1(\theRegs/completionDataOut[3][41] ), .A2(n3474), .B1(
        \theRegs/completionDataOut[1][41] ), .B2(n3446), .ZN(n2966) );
  AOI22D2 U3241 ( .A1(\theRegs/completionDataOut[7][1] ), .A2(n3346), .B1(
        \theRegs/completionDataOut[4][1] ), .B2(n3523), .ZN(n3124) );
  AOI22D2 U3954 ( .A1(\theRegs/completionDataOut[3][32] ), .A2(n3398), .B1(
        \theRegs/completionDataOut[1][32] ), .B2(n3379), .ZN(n3002) );
  AOI22D2 U4034 ( .A1(\theRegs/completionDataOut[3][47] ), .A2(n3558), .B1(
        \theRegs/completionDataOut[1][47] ), .B2(n3521), .ZN(n2942) );
  AOI22D2 U3682 ( .A1(\theRegs/completionDataOut[7][42] ), .A2(n3274), .B1(
        \theRegs/completionDataOut[6][42] ), .B2(n3268), .ZN(n2687) );
  AOI22D2 U4027 ( .A1(\theRegs/completionDataOut[7][46] ), .A2(n3282), .B1(
        \theRegs/completionDataOut[4][46] ), .B2(n3270), .ZN(n2944) );
  AOI22D2 U4077 ( .A1(\theRegs/completionDataOut[7][56] ), .A2(n3282), .B1(
        \theRegs/completionDataOut[4][56] ), .B2(n3270), .ZN(n2904) );
  AOI22D2 U3664 ( .A1(\theRegs/completionDataOut[3][46] ), .A2(n3458), .B1(
        \theRegs/completionDataOut[1][46] ), .B2(n3526), .ZN(n2673) );
  AOI22D2 U3729 ( .A1(\theRegs/completionDataOut[3][55] ), .A2(n3485), .B1(
        \theRegs/completionDataOut[1][55] ), .B2(n3557), .ZN(n2637) );
  AOI22D2 U3153 ( .A1(\theRegs/completionDataOut[3][19] ), .A2(n3398), .B1(
        \theRegs/completionDataOut[1][19] ), .B2(n3379), .ZN(n3054) );
  AOI22D2 U3862 ( .A1(\theRegs/completionDataOut[7][19] ), .A2(n3455), .B1(
        \theRegs/completionDataOut[6][19] ), .B2(n3487), .ZN(n2779) );
  AOI22D2 U3792 ( .A1(\theRegs/completionDataOut[7][33] ), .A2(n3455), .B1(
        \theRegs/completionDataOut[6][33] ), .B2(n3487), .ZN(n2723) );
  AOI22D2 U3654 ( .A1(\theRegs/completionDataOut[3][48] ), .A2(n3485), .B1(
        \theRegs/completionDataOut[1][48] ), .B2(n3557), .ZN(n2665) );
  AOI22D2 U3236 ( .A1(\theRegs/completionDataOut[7][2] ), .A2(n3347), .B1(
        \theRegs/completionDataOut[4][2] ), .B2(n3540), .ZN(n3120) );
  AOI22D2 U4002 ( .A1(\theRegs/completionDataOut[7][41] ), .A2(n3282), .B1(
        \theRegs/completionDataOut[4][41] ), .B2(n3270), .ZN(n2964) );
  AOI22D2 U3595 ( .A1(n3345), .A2(\theRegs/completionDataOut[4][11] ), .B1(
        n3356), .B2(\theRegs/completionDataOut[0][11] ), .ZN(n2354) );
  AOI22D2 U3819 ( .A1(\theRegs/completionDataOut[3][28] ), .A2(n3437), .B1(
        \theRegs/completionDataOut[1][28] ), .B2(n3406), .ZN(n2745) );
  AOI22D2 U4039 ( .A1(\theRegs/completionDataOut[3][48] ), .A2(n3558), .B1(
        \theRegs/completionDataOut[1][48] ), .B2(n3521), .ZN(n2938) );
  AOI22D2 U4079 ( .A1(\theRegs/completionDataOut[3][56] ), .A2(n3558), .B1(
        \theRegs/completionDataOut[1][56] ), .B2(n3521), .ZN(n2906) );
  AOI22D2 U3912 ( .A1(\theRegs/completionDataOut[7][9] ), .A2(n3455), .B1(
        \theRegs/completionDataOut[6][9] ), .B2(n3487), .ZN(n2819) );
  AOI22D2 U4074 ( .A1(\theRegs/completionDataOut[3][55] ), .A2(n3558), .B1(
        \theRegs/completionDataOut[1][55] ), .B2(n3521), .ZN(n2910) );
  AOI22D2 U4152 ( .A1(\theRegs/completionDataOut[3][59] ), .A2(n3585), .B1(
        \theRegs/completionDataOut[1][59] ), .B2(n3543), .ZN(n2894) );
  AOI22D2 U3659 ( .A1(\theRegs/completionDataOut[3][47] ), .A2(n3485), .B1(
        \theRegs/completionDataOut[1][47] ), .B2(n3557), .ZN(n2669) );
  AOI22D2 U3151 ( .A1(\theRegs/completionDataOut[7][19] ), .A2(n3347), .B1(
        \theRegs/completionDataOut[4][19] ), .B2(n3540), .ZN(n3052) );
  AOI22D2 U4084 ( .A1(\theRegs/completionDataOut[3][57] ), .A2(n3585), .B1(
        \theRegs/completionDataOut[1][57] ), .B2(n3543), .ZN(n2902) );
  AOI22D2 U3754 ( .A1(\theRegs/completionDataOut[3][49] ), .A2(n3485), .B1(
        \theRegs/completionDataOut[1][49] ), .B2(n3557), .ZN(n2661) );
  AOI22D2 U3198 ( .A1(\theRegs/completionDataOut[3][10] ), .A2(n3398), .B1(
        \theRegs/completionDataOut[1][10] ), .B2(n3379), .ZN(n3090) );
  AOI22D2 U3490 ( .A1(n3345), .A2(\theRegs/completionDataOut[4][32] ), .B1(
        n3385), .B2(\theRegs/completionDataOut[0][32] ), .ZN(n2438) );
  AOI22D2 U3724 ( .A1(\theRegs/completionDataOut[3][54] ), .A2(n3485), .B1(
        \theRegs/completionDataOut[1][54] ), .B2(n3557), .ZN(n2641) );
  AOI22D2 U3739 ( .A1(\theRegs/completionDataOut[3][57] ), .A2(n3542), .B1(
        \theRegs/completionDataOut[1][57] ), .B2(n3584), .ZN(n2629) );
  AOI22D2 U3166 ( .A1(\theRegs/completionDataOut[7][16] ), .A2(n3347), .B1(
        \theRegs/completionDataOut[4][16] ), .B2(n3540), .ZN(n3064) );
  AOI22D2 U3432 ( .A1(n3363), .A2(\theRegs/completionDataOut[6][43] ), .B1(
        n3304), .B2(\theRegs/completionDataOut[7][43] ), .ZN(n2479) );
  AOI22D2 U3649 ( .A1(\theRegs/completionDataOut[3][63] ), .A2(n3542), .B1(
        \theRegs/completionDataOut[1][63] ), .B2(n3584), .ZN(n2605) );
  CKBD4 U4196 ( .I(n2178), .Z(n3316) );
  AOI22D2 U3662 ( .A1(\theRegs/completionDataOut[7][46] ), .A2(n3274), .B1(
        \theRegs/completionDataOut[6][46] ), .B2(n3268), .ZN(n2671) );
  AOI22D2 U3727 ( .A1(\theRegs/completionDataOut[7][55] ), .A2(n3274), .B1(
        \theRegs/completionDataOut[6][55] ), .B2(n3268), .ZN(n2635) );
  AOI22D2 U3359 ( .A1(\theRegs/completionDataOut[3][28] ), .A2(n3398), .B1(
        \theRegs/completionDataOut[1][28] ), .B2(n3379), .ZN(n3018) );
  AOI22D2 U3437 ( .A1(n3363), .A2(\theRegs/completionDataOut[6][42] ), .B1(
        n3625), .B2(\theRegs/completionDataOut[7][42] ), .ZN(n2475) );
  CKBD3 U4216 ( .I(n2182), .Z(n3326) );
  AOI22D2 U3417 ( .A1(n3363), .A2(\theRegs/completionDataOut[6][46] ), .B1(
        n3625), .B2(\theRegs/completionDataOut[7][46] ), .ZN(n2491) );
  AOI22D2 U3957 ( .A1(\theRegs/completionDataOut[7][33] ), .A2(n3347), .B1(
        \theRegs/completionDataOut[4][33] ), .B2(n3540), .ZN(n2996) );
  AOI22D2 U3834 ( .A1(\theRegs/completionDataOut[3][25] ), .A2(n3561), .B1(
        \theRegs/completionDataOut[1][25] ), .B2(n3488), .ZN(n2757) );
  AOI22D2 U3807 ( .A1(\theRegs/completionDataOut[7][30] ), .A2(n3455), .B1(
        \theRegs/completionDataOut[6][30] ), .B2(n3487), .ZN(n2735) );
  AOI22D2 U3213 ( .A1(\theRegs/completionDataOut[3][7] ), .A2(n3398), .B1(
        \theRegs/completionDataOut[1][7] ), .B2(n3379), .ZN(n3102) );
  AOI22D2 U3962 ( .A1(\theRegs/completionDataOut[7][34] ), .A2(n3347), .B1(
        \theRegs/completionDataOut[4][34] ), .B2(n3540), .ZN(n2992) );
  AOI22D2 U3997 ( .A1(\theRegs/completionDataOut[7][40] ), .A2(n3447), .B1(
        \theRegs/completionDataOut[4][40] ), .B2(n3415), .ZN(n2968) );
  BUFFD2 U4192 ( .I(n2181), .Z(n3314) );
  AOI22D2 U4044 ( .A1(\theRegs/completionDataOut[3][49] ), .A2(n3585), .B1(
        \theRegs/completionDataOut[1][49] ), .B2(n3543), .ZN(n2934) );
  AOI22D2 U3515 ( .A1(n3345), .A2(\theRegs/completionDataOut[4][27] ), .B1(
        n3385), .B2(\theRegs/completionDataOut[0][27] ), .ZN(n2418) );
  AOI22D2 U4097 ( .A1(\theRegs/completionDataOut[7][64] ), .A2(n3447), .B1(
        \theRegs/completionDataOut[4][64] ), .B2(n3415), .ZN(n2872) );
  AOI22D2 U3872 ( .A1(\theRegs/completionDataOut[7][17] ), .A2(n3455), .B1(
        \theRegs/completionDataOut[6][17] ), .B2(n3487), .ZN(n2787) );
  AOI22D2 U3211 ( .A1(\theRegs/completionDataOut[7][7] ), .A2(n3353), .B1(
        \theRegs/completionDataOut[4][7] ), .B2(n3592), .ZN(n3100) );
  AOI221D4 U4848 ( .A1(n3793), .A2(tail[0]), .B1(n3312), .B2(n3238), .C(n2264), 
        .ZN(n1402) );
  AOI22D2 U4150 ( .A1(\theRegs/completionDataOut[7][59] ), .A2(n3447), .B1(
        \theRegs/completionDataOut[4][59] ), .B2(n3415), .ZN(n2892) );
  AOI22D2 U3442 ( .A1(n3363), .A2(\theRegs/completionDataOut[6][41] ), .B1(
        n3625), .B2(\theRegs/completionDataOut[7][41] ), .ZN(n2471) );
  AOI22D2 U3769 ( .A1(\theRegs/completionDataOut[3][38] ), .A2(n3542), .B1(
        \theRegs/completionDataOut[1][38] ), .B2(n3584), .ZN(n2705) );
  AOI22D2 U3176 ( .A1(\theRegs/completionDataOut[7][14] ), .A2(n3353), .B1(
        \theRegs/completionDataOut[4][14] ), .B2(n3592), .ZN(n3072) );
  AOI22D2 U4069 ( .A1(\theRegs/completionDataOut[3][54] ), .A2(n3585), .B1(
        \theRegs/completionDataOut[1][54] ), .B2(n3543), .ZN(n2914) );
  AOI22D2 U3123 ( .A1(\theRegs/completionDataOut[3][25] ), .A2(n3424), .B1(
        \theRegs/completionDataOut[1][25] ), .B2(n3454), .ZN(n3030) );
  AOI22D2 U3677 ( .A1(\theRegs/completionDataOut[7][43] ), .A2(n3274), .B1(
        \theRegs/completionDataOut[6][43] ), .B2(n3407), .ZN(n2683) );
  AOI22D2 U3226 ( .A1(\theRegs/completionDataOut[7][4] ), .A2(n3353), .B1(
        \theRegs/completionDataOut[4][4] ), .B2(n3592), .ZN(n3112) );
  CKBD3 U4219 ( .I(n2187), .Z(n3329) );
  AOI22D2 U4082 ( .A1(\theRegs/completionDataOut[7][57] ), .A2(n3447), .B1(
        \theRegs/completionDataOut[4][57] ), .B2(n3415), .ZN(n2900) );
  AOI22D2 U3667 ( .A1(\theRegs/completionDataOut[7][45] ), .A2(n3459), .B1(
        \theRegs/completionDataOut[6][45] ), .B2(n3407), .ZN(n2675) );
  CKBD3 U4227 ( .I(n2184), .Z(n3337) );
  AOI22D2 U3427 ( .A1(n3363), .A2(\theRegs/completionDataOut[6][44] ), .B1(
        n3625), .B2(\theRegs/completionDataOut[7][44] ), .ZN(n2483) );
  AOI22D2 U3869 ( .A1(\theRegs/completionDataOut[3][18] ), .A2(n3561), .B1(
        \theRegs/completionDataOut[1][18] ), .B2(n3488), .ZN(n2785) );
  AOI22D2 U3645 ( .A1(n3298), .A2(\theRegs/completionDataOut[4][1] ), .B1(
        n3422), .B2(\theRegs/completionDataOut[0][1] ), .ZN(n2314) );
  AOI22D2 U3188 ( .A1(\theRegs/completionDataOut[3][12] ), .A2(n3424), .B1(
        \theRegs/completionDataOut[1][12] ), .B2(n3454), .ZN(n3082) );
  AOI22D2 U3732 ( .A1(\theRegs/completionDataOut[7][56] ), .A2(n3459), .B1(
        \theRegs/completionDataOut[6][56] ), .B2(n3490), .ZN(n2631) );
  AOI22D2 U3191 ( .A1(\theRegs/completionDataOut[7][11] ), .A2(n3358), .B1(
        \theRegs/completionDataOut[4][11] ), .B2(n3658), .ZN(n3084) );
  AOI22D2 U3555 ( .A1(n3345), .A2(\theRegs/completionDataOut[4][19] ), .B1(
        n3422), .B2(\theRegs/completionDataOut[0][19] ), .ZN(n2386) );
  AOI22D2 U3694 ( .A1(\theRegs/completionDataOut[3][40] ), .A2(n3542), .B1(
        \theRegs/completionDataOut[1][40] ), .B2(n3584), .ZN(n2697) );
  AOI22D2 U3171 ( .A1(\theRegs/completionDataOut[7][15] ), .A2(n3358), .B1(
        \theRegs/completionDataOut[4][15] ), .B2(n3658), .ZN(n3068) );
  AOI22D2 U4124 ( .A1(\theRegs/completionDataOut[3][60] ), .A2(n3630), .B1(
        \theRegs/completionDataOut[1][60] ), .B2(n3674), .ZN(n2617) );
  AOI22D2 U3672 ( .A1(\theRegs/completionDataOut[7][44] ), .A2(n3459), .B1(
        \theRegs/completionDataOut[6][44] ), .B2(n3490), .ZN(n2679) );
  AOI22D2 U3924 ( .A1(\theRegs/completionDataOut[3][7] ), .A2(n3598), .B1(
        \theRegs/completionDataOut[1][7] ), .B2(n3519), .ZN(n2829) );
  AOI22D2 U4007 ( .A1(\theRegs/completionDataOut[7][29] ), .A2(n3358), .B1(
        \theRegs/completionDataOut[4][29] ), .B2(n3658), .ZN(n3012) );
  AOI22D2 U3932 ( .A1(\theRegs/completionDataOut[7][5] ), .A2(n3463), .B1(
        \theRegs/completionDataOut[6][5] ), .B2(n3497), .ZN(n2835) );
  AOI22D2 U3372 ( .A1(n3370), .A2(\theRegs/completionDataOut[6][55] ), .B1(
        n3625), .B2(\theRegs/completionDataOut[7][55] ), .ZN(n2527) );
  AOI22D2 U3181 ( .A1(\theRegs/completionDataOut[7][13] ), .A2(n3358), .B1(
        \theRegs/completionDataOut[4][13] ), .B2(n3658), .ZN(n3076) );
  AOI22D2 U3999 ( .A1(\theRegs/completionDataOut[3][40] ), .A2(n3675), .B1(
        \theRegs/completionDataOut[1][40] ), .B2(n3631), .ZN(n2970) );
  AOI22D2 U3592 ( .A1(n3457), .A2(\theRegs/completionDataOut[6][11] ), .B1(
        n3642), .B2(\theRegs/completionDataOut[7][11] ), .ZN(n2351) );
  AOI22D2 U3722 ( .A1(\theRegs/completionDataOut[7][54] ), .A2(n3459), .B1(
        \theRegs/completionDataOut[6][54] ), .B2(n3490), .ZN(n2639) );
  AOI22D2 U4104 ( .A1(\theRegs/completionDataOut[3][0] ), .A2(n3598), .B1(
        \theRegs/completionDataOut[1][0] ), .B2(n3519), .ZN(n2865) );
  AOI22D2 U4092 ( .A1(\theRegs/completionDataOut[7][58] ), .A2(n3469), .B1(
        \theRegs/completionDataOut[4][58] ), .B2(n3444), .ZN(n2896) );
  AOI22D2 U3163 ( .A1(\theRegs/completionDataOut[3][17] ), .A2(n3424), .B1(
        \theRegs/completionDataOut[1][17] ), .B2(n3454), .ZN(n3062) );
  AOI22D2 U3362 ( .A1(n3370), .A2(\theRegs/completionDataOut[6][57] ), .B1(
        n3661), .B2(\theRegs/completionDataOut[7][57] ), .ZN(n2535) );
  AOI22D2 U3575 ( .A1(n3345), .A2(\theRegs/completionDataOut[4][15] ), .B1(
        n3422), .B2(\theRegs/completionDataOut[0][15] ), .ZN(n2370) );
  AOI22D2 U3692 ( .A1(\theRegs/completionDataOut[7][40] ), .A2(n3459), .B1(
        \theRegs/completionDataOut[6][40] ), .B2(n3490), .ZN(n2695) );
  AOI22D2 U3897 ( .A1(\theRegs/completionDataOut[7][12] ), .A2(n3463), .B1(
        \theRegs/completionDataOut[6][12] ), .B2(n3497), .ZN(n2807) );
  AOI22D2 U3922 ( .A1(\theRegs/completionDataOut[7][7] ), .A2(n3463), .B1(
        \theRegs/completionDataOut[6][7] ), .B2(n3497), .ZN(n2827) );
  AOI22D2 U3570 ( .A1(n3348), .A2(\theRegs/completionDataOut[4][16] ), .B1(
        n3422), .B2(\theRegs/completionDataOut[0][16] ), .ZN(n2374) );
  AOI22D2 U3714 ( .A1(\theRegs/completionDataOut[3][52] ), .A2(n3630), .B1(
        \theRegs/completionDataOut[1][52] ), .B2(n3674), .ZN(n2649) );
  AOI22D2 U3735 ( .A1(\theRegs/completionDataOut[2][56] ), .A2(n3279), .B1(
        \theRegs/completionDataOut[0][56] ), .B2(n3263), .ZN(n2634) );
  AOI22D2 U3707 ( .A1(\theRegs/completionDataOut[7][51] ), .A2(n3465), .B1(
        \theRegs/completionDataOut[6][51] ), .B2(n3502), .ZN(n2651) );
  AOI22D2 U3186 ( .A1(\theRegs/completionDataOut[7][12] ), .A2(n3358), .B1(
        \theRegs/completionDataOut[4][12] ), .B2(n3658), .ZN(n3080) );
  AOI22D2 U4087 ( .A1(\theRegs/completionDataOut[7][42] ), .A2(n3469), .B1(
        \theRegs/completionDataOut[4][42] ), .B2(n3444), .ZN(n2960) );
  AO21D2 U2270 ( .A1(n3140), .A2(n3298), .B(reset_i), .Z(n2223) );
  AOI22D2 U3505 ( .A1(n3354), .A2(\theRegs/completionDataOut[4][29] ), .B1(
        n3422), .B2(\theRegs/completionDataOut[0][29] ), .ZN(n2426) );
  AOI22D2 U4145 ( .A1(\theRegs/completionDataOut[7][61] ), .A2(n3469), .B1(
        \theRegs/completionDataOut[4][61] ), .B2(n3444), .ZN(n2884) );
  CKBD3 U4231 ( .I(n2188), .Z(n3341) );
  AOI22D2 U3909 ( .A1(\theRegs/completionDataOut[3][10] ), .A2(n3598), .B1(
        \theRegs/completionDataOut[1][10] ), .B2(n3519), .ZN(n2817) );
  AOI22D2 U3882 ( .A1(\theRegs/completionDataOut[7][15] ), .A2(n3463), .B1(
        \theRegs/completionDataOut[6][15] ), .B2(n3497), .ZN(n2795) );
  AOI22D2 U3744 ( .A1(\theRegs/completionDataOut[3][58] ), .A2(n3630), .B1(
        \theRegs/completionDataOut[1][58] ), .B2(n3674), .ZN(n2625) );
  AOI22D2 U3719 ( .A1(\theRegs/completionDataOut[3][53] ), .A2(n3630), .B1(
        \theRegs/completionDataOut[1][53] ), .B2(n3674), .ZN(n2645) );
  AOI22D2 U3702 ( .A1(\theRegs/completionDataOut[7][50] ), .A2(n3465), .B1(
        \theRegs/completionDataOut[6][50] ), .B2(n3502), .ZN(n2655) );
  AOI22D2 U3367 ( .A1(n3370), .A2(\theRegs/completionDataOut[6][56] ), .B1(
        n3661), .B2(\theRegs/completionDataOut[7][56] ), .ZN(n2531) );
  CKBD3 U4212 ( .I(n2185), .Z(n3322) );
  AOI22D2 U3246 ( .A1(\theRegs/completionDataOut[7][0] ), .A2(n3368), .B1(
        \theRegs/completionDataOut[4][0] ), .B2(n3714), .ZN(n3136) );
  AOI22D2 U3231 ( .A1(\theRegs/completionDataOut[7][3] ), .A2(n3368), .B1(
        \theRegs/completionDataOut[4][3] ), .B2(n3714), .ZN(n3116) );
  AOI22D2 U3248 ( .A1(\theRegs/completionDataOut[3][0] ), .A2(n3424), .B1(
        \theRegs/completionDataOut[1][0] ), .B2(n3454), .ZN(n3138) );
  AOI22D2 U3904 ( .A1(\theRegs/completionDataOut[3][11] ), .A2(n3598), .B1(
        \theRegs/completionDataOut[1][11] ), .B2(n3519), .ZN(n2813) );
  AOI22D2 U3158 ( .A1(\theRegs/completionDataOut[3][18] ), .A2(n3424), .B1(
        \theRegs/completionDataOut[1][18] ), .B2(n3454), .ZN(n3058) );
  AOI22D2 U4059 ( .A1(\theRegs/completionDataOut[3][52] ), .A2(n3675), .B1(
        \theRegs/completionDataOut[1][52] ), .B2(n3631), .ZN(n2922) );
  AOI22D2 U3510 ( .A1(n3354), .A2(\theRegs/completionDataOut[4][28] ), .B1(
        n3432), .B2(\theRegs/completionDataOut[0][28] ), .ZN(n2422) );
  AOI22D2 U3877 ( .A1(\theRegs/completionDataOut[7][16] ), .A2(n3463), .B1(
        \theRegs/completionDataOut[6][16] ), .B2(n3497), .ZN(n2791) );
  AOI22D2 U4017 ( .A1(\theRegs/completionDataOut[7][44] ), .A2(n3469), .B1(
        \theRegs/completionDataOut[4][44] ), .B2(n3444), .ZN(n2952) );
  BUFFD1 U4217 ( .I(n4115), .Z(n3327) );
  AOI22D2 U3992 ( .A1(\theRegs/completionDataOut[7][39] ), .A2(n3553), .B1(
        \theRegs/completionDataOut[4][39] ), .B2(n3518), .ZN(n2972) );
  AOI22D2 U3884 ( .A1(\theRegs/completionDataOut[3][15] ), .A2(n3598), .B1(
        \theRegs/completionDataOut[1][15] ), .B2(n3519), .ZN(n2797) );
  AOI22D2 U3892 ( .A1(\theRegs/completionDataOut[7][13] ), .A2(n3550), .B1(
        \theRegs/completionDataOut[6][13] ), .B2(n3594), .ZN(n2803) );
  AOI22D2 U3687 ( .A1(\theRegs/completionDataOut[7][41] ), .A2(n3465), .B1(
        \theRegs/completionDataOut[6][41] ), .B2(n3502), .ZN(n2691) );
  AOI22D2 U4130 ( .A1(\theRegs/completionDataOut[7][62] ), .A2(n3553), .B1(
        \theRegs/completionDataOut[4][62] ), .B2(n3518), .ZN(n2880) );
  AOI22D2 U3412 ( .A1(n3370), .A2(\theRegs/completionDataOut[6][47] ), .B1(
        n3661), .B2(\theRegs/completionDataOut[7][47] ), .ZN(n2495) );
  AOI22D2 U3173 ( .A1(\theRegs/completionDataOut[3][15] ), .A2(n3435), .B1(
        \theRegs/completionDataOut[1][15] ), .B2(n3467), .ZN(n3070) );
  AOI22D2 U3937 ( .A1(\theRegs/completionDataOut[7][4] ), .A2(n3581), .B1(
        \theRegs/completionDataOut[6][4] ), .B2(n3618), .ZN(n2839) );
  AOI22D2 U4012 ( .A1(\theRegs/completionDataOut[7][43] ), .A2(n3553), .B1(
        \theRegs/completionDataOut[4][43] ), .B2(n3518), .ZN(n2956) );
  AOI22D2 U3902 ( .A1(\theRegs/completionDataOut[7][11] ), .A2(n3581), .B1(
        \theRegs/completionDataOut[6][11] ), .B2(n3618), .ZN(n2811) );
  AOI22D2 U3565 ( .A1(n3354), .A2(\theRegs/completionDataOut[4][17] ), .B1(
        n3432), .B2(\theRegs/completionDataOut[0][17] ), .ZN(n2378) );
  AOI22D2 U3742 ( .A1(\theRegs/completionDataOut[7][58] ), .A2(n3465), .B1(
        \theRegs/completionDataOut[6][58] ), .B2(n3502), .ZN(n2623) );
  CKBD4 U4228 ( .I(n2184), .Z(n3338) );
  AOI22D2 U3887 ( .A1(\theRegs/completionDataOut[7][14] ), .A2(n3581), .B1(
        \theRegs/completionDataOut[6][14] ), .B2(n3618), .ZN(n2799) );
  AOI22D2 U3350 ( .A1(n3298), .A2(\theRegs/completionDataOut[4][59] ), .B1(
        n3275), .B2(\theRegs/completionDataOut[0][59] ), .ZN(n2546) );
  AOI22D2 U3168 ( .A1(\theRegs/completionDataOut[3][16] ), .A2(n3435), .B1(
        \theRegs/completionDataOut[1][16] ), .B2(n3467), .ZN(n3066) );
  AOI22D2 U3889 ( .A1(\theRegs/completionDataOut[3][14] ), .A2(n3619), .B1(
        \theRegs/completionDataOut[1][14] ), .B2(n3582), .ZN(n2801) );
  AOI22D2 U3657 ( .A1(\theRegs/completionDataOut[7][47] ), .A2(n3554), .B1(
        \theRegs/completionDataOut[6][47] ), .B2(n3596), .ZN(n2667) );
  AOI22D2 U4119 ( .A1(\theRegs/completionDataOut[3][3] ), .A2(n3619), .B1(
        \theRegs/completionDataOut[1][3] ), .B2(n3582), .ZN(n2845) );
  AOI22D2 U4135 ( .A1(\theRegs/completionDataOut[7][63] ), .A2(n3553), .B1(
        \theRegs/completionDataOut[4][63] ), .B2(n3518), .ZN(n2876) );
  AOI22D2 U3335 ( .A1(n3609), .A2(\theRegs/completionDataOut[4][62] ), .B1(
        n3275), .B2(\theRegs/completionDataOut[0][62] ), .ZN(n2558) );
  AOI22D2 U4140 ( .A1(\theRegs/completionDataOut[7][60] ), .A2(n3570), .B1(
        \theRegs/completionDataOut[4][60] ), .B2(n3532), .ZN(n2888) );
  AOI22D2 U3233 ( .A1(\theRegs/completionDataOut[3][3] ), .A2(n3435), .B1(
        \theRegs/completionDataOut[1][3] ), .B2(n3467), .ZN(n3118) );
  AOI22D2 U3445 ( .A1(n3609), .A2(\theRegs/completionDataOut[4][41] ), .B1(
        n3275), .B2(\theRegs/completionDataOut[0][41] ), .ZN(n2474) );
  AOI22D2 U3927 ( .A1(\theRegs/completionDataOut[7][6] ), .A2(n3581), .B1(
        \theRegs/completionDataOut[6][6] ), .B2(n3618), .ZN(n2831) );
  AOI22D2 U3567 ( .A1(n3457), .A2(\theRegs/completionDataOut[6][16] ), .B1(
        n3642), .B2(\theRegs/completionDataOut[7][16] ), .ZN(n2371) );
  AOI22D2 U4032 ( .A1(\theRegs/completionDataOut[7][47] ), .A2(n3570), .B1(
        \theRegs/completionDataOut[4][47] ), .B2(n3532), .ZN(n2940) );
  AOI22D2 U3967 ( .A1(\theRegs/completionDataOut[7][35] ), .A2(n3570), .B1(
        \theRegs/completionDataOut[4][35] ), .B2(n3532), .ZN(n2988) );
  AOI22D2 U3347 ( .A1(n3370), .A2(\theRegs/completionDataOut[6][59] ), .B1(
        n3661), .B2(\theRegs/completionDataOut[7][59] ), .ZN(n2543) );
  AOI22D2 U3297 ( .A1(n3377), .A2(\theRegs/completionDataOut[6][69] ), .B1(
        n3661), .B2(\theRegs/completionDataOut[7][69] ), .ZN(n2590) );
  AOI22D2 U4054 ( .A1(\theRegs/completionDataOut[3][51] ), .A2(n3675), .B1(
        \theRegs/completionDataOut[1][51] ), .B2(n3631), .ZN(n2926) );
  AOI22D2 U3325 ( .A1(n3609), .A2(\theRegs/completionDataOut[4][64] ), .B1(
        n3275), .B2(\theRegs/completionDataOut[0][64] ), .ZN(n2566) );
  AOI22D2 U3709 ( .A1(\theRegs/completionDataOut[3][51] ), .A2(n3650), .B1(
        \theRegs/completionDataOut[1][51] ), .B2(n3692), .ZN(n2653) );
  AOI22D2 U3370 ( .A1(n3354), .A2(\theRegs/completionDataOut[4][56] ), .B1(
        n3411), .B2(\theRegs/completionDataOut[0][56] ), .ZN(n2534) );
  AOI22D2 U3894 ( .A1(\theRegs/completionDataOut[3][13] ), .A2(n3619), .B1(
        \theRegs/completionDataOut[1][13] ), .B2(n3582), .ZN(n2805) );
  AOI22D2 U3737 ( .A1(\theRegs/completionDataOut[7][57] ), .A2(n3554), .B1(
        \theRegs/completionDataOut[6][57] ), .B2(n3596), .ZN(n2627) );
  AOI22D2 U3377 ( .A1(n3377), .A2(\theRegs/completionDataOut[6][54] ), .B1(
        n3724), .B2(\theRegs/completionDataOut[7][54] ), .ZN(n2523) );
  AOI22D2 U4064 ( .A1(\theRegs/completionDataOut[3][53] ), .A2(n3675), .B1(
        \theRegs/completionDataOut[1][53] ), .B2(n3631), .ZN(n2918) );
  AOI22D2 U3577 ( .A1(n3457), .A2(\theRegs/completionDataOut[6][14] ), .B1(
        n3642), .B2(\theRegs/completionDataOut[7][14] ), .ZN(n2363) );
  AOI22D2 U3560 ( .A1(n3354), .A2(\theRegs/completionDataOut[4][18] ), .B1(
        n3432), .B2(\theRegs/completionDataOut[0][18] ), .ZN(n2382) );
  CKND2 U2478 ( .I(n3212), .ZN(n3213) );
  AOI22D2 U3562 ( .A1(n3457), .A2(\theRegs/completionDataOut[6][17] ), .B1(
        n3656), .B2(\theRegs/completionDataOut[7][17] ), .ZN(n2375) );
  AOI22D2 U3397 ( .A1(n3377), .A2(\theRegs/completionDataOut[6][50] ), .B1(
        n3724), .B2(\theRegs/completionDataOut[7][50] ), .ZN(n2507) );
  AOI22D2 U3770 ( .A1(\theRegs/completionDataOut[2][38] ), .A2(n3280), .B1(
        \theRegs/completionDataOut[0][38] ), .B2(n3264), .ZN(n2706) );
  AOI22D2 U3422 ( .A1(n3377), .A2(\theRegs/completionDataOut[6][45] ), .B1(
        n3724), .B2(\theRegs/completionDataOut[7][45] ), .ZN(n2487) );
  AOI22D2 U3475 ( .A1(n3609), .A2(\theRegs/completionDataOut[4][35] ), .B1(
        n3411), .B2(\theRegs/completionDataOut[0][35] ), .ZN(n2450) );
  AOI22D2 U3899 ( .A1(\theRegs/completionDataOut[3][12] ), .A2(n3619), .B1(
        \theRegs/completionDataOut[1][12] ), .B2(n3582), .ZN(n2809) );
  AOI22D2 U3178 ( .A1(\theRegs/completionDataOut[3][14] ), .A2(n3435), .B1(
        \theRegs/completionDataOut[1][14] ), .B2(n3467), .ZN(n3074) );
  AOI22D2 U3447 ( .A1(n3400), .A2(\theRegs/completionDataOut[6][40] ), .B1(
        n3724), .B2(\theRegs/completionDataOut[7][40] ), .ZN(n2467) );
  AOI22D2 U3352 ( .A1(n3400), .A2(\theRegs/completionDataOut[6][58] ), .B1(
        n3754), .B2(\theRegs/completionDataOut[7][58] ), .ZN(n2539) );
  AOI22D2 U3435 ( .A1(n3733), .A2(\theRegs/completionDataOut[4][43] ), .B1(
        n3411), .B2(\theRegs/completionDataOut[0][43] ), .ZN(n2482) );
  AOI22D2 U3772 ( .A1(\theRegs/completionDataOut[7][37] ), .A2(n3554), .B1(
        \theRegs/completionDataOut[6][37] ), .B2(n3596), .ZN(n2707) );
  AOI22D2 U3403 ( .A1(n3301), .A2(\theRegs/completionDataOut[5][49] ), .B1(
        n3288), .B2(\theRegs/completionDataOut[3][49] ), .ZN(n2504) );
  AOI22D2 U3580 ( .A1(n3359), .A2(\theRegs/completionDataOut[4][14] ), .B1(
        n3432), .B2(\theRegs/completionDataOut[0][14] ), .ZN(n2366) );
  AOI22D2 U3630 ( .A1(n3733), .A2(\theRegs/completionDataOut[4][4] ), .B1(
        n3482), .B2(\theRegs/completionDataOut[0][4] ), .ZN(n2326) );
  INR2XD2 U3082 ( .A1(n2233), .B1(n2232), .ZN(n2234) );
  AOI22D2 U3183 ( .A1(\theRegs/completionDataOut[3][13] ), .A2(n3435), .B1(
        \theRegs/completionDataOut[1][13] ), .B2(n3467), .ZN(n3078) );
  AOI22D2 U3879 ( .A1(\theRegs/completionDataOut[3][16] ), .A2(n3619), .B1(
        \theRegs/completionDataOut[1][16] ), .B2(n3582), .ZN(n2793) );
  AOI22D2 U3458 ( .A1(n3352), .A2(\theRegs/completionDataOut[5][38] ), .B1(
        n3286), .B2(\theRegs/completionDataOut[3][38] ), .ZN(n2460) );
  AOI22D2 U3587 ( .A1(n3494), .A2(\theRegs/completionDataOut[6][12] ), .B1(
        n3656), .B2(\theRegs/completionDataOut[7][12] ), .ZN(n2355) );
  AOI22D2 U3557 ( .A1(n3494), .A2(\theRegs/completionDataOut[6][18] ), .B1(
        n3656), .B2(\theRegs/completionDataOut[7][18] ), .ZN(n2379) );
  CKBD3 U4213 ( .I(n2185), .Z(n3323) );
  AOI22D2 U3193 ( .A1(\theRegs/completionDataOut[3][11] ), .A2(n3549), .B1(
        \theRegs/completionDataOut[1][11] ), .B2(n3514), .ZN(n3086) );
  AOI22D2 U3330 ( .A1(n3771), .A2(\theRegs/completionDataOut[4][63] ), .B1(
        n3456), .B2(\theRegs/completionDataOut[0][63] ), .ZN(n2562) );
  AOI22D2 U3552 ( .A1(n3494), .A2(\theRegs/completionDataOut[6][19] ), .B1(
        n3656), .B2(\theRegs/completionDataOut[7][19] ), .ZN(n2383) );
  AOI22D2 U3602 ( .A1(n3374), .A2(\theRegs/completionDataOut[6][9] ), .B1(
        n3656), .B2(\theRegs/completionDataOut[7][9] ), .ZN(n2343) );
  AOI22D2 U3477 ( .A1(n3400), .A2(\theRegs/completionDataOut[6][34] ), .B1(
        n3754), .B2(\theRegs/completionDataOut[7][34] ), .ZN(n2443) );
  AOI22D2 U3440 ( .A1(n3771), .A2(\theRegs/completionDataOut[4][42] ), .B1(
        n3456), .B2(\theRegs/completionDataOut[0][42] ), .ZN(n2478) );
  AOI22D2 U3582 ( .A1(n3494), .A2(\theRegs/completionDataOut[6][13] ), .B1(
        n3656), .B2(\theRegs/completionDataOut[7][13] ), .ZN(n2359) );
  AOI22D2 U3640 ( .A1(n3771), .A2(\theRegs/completionDataOut[4][2] ), .B1(
        n3482), .B2(\theRegs/completionDataOut[0][2] ), .ZN(n2318) );
  AOI22D2 U3368 ( .A1(n3301), .A2(\theRegs/completionDataOut[5][56] ), .B1(
        n3288), .B2(\theRegs/completionDataOut[3][56] ), .ZN(n2532) );
  AOI22D2 U3572 ( .A1(n3494), .A2(\theRegs/completionDataOut[6][15] ), .B1(
        n3725), .B2(\theRegs/completionDataOut[7][15] ), .ZN(n2367) );
  AOI22D2 U3355 ( .A1(n3359), .A2(\theRegs/completionDataOut[4][58] ), .B1(
        n3456), .B2(\theRegs/completionDataOut[0][58] ), .ZN(n2542) );
  AOI22D2 U3340 ( .A1(n3771), .A2(\theRegs/completionDataOut[4][61] ), .B1(
        n3456), .B2(\theRegs/completionDataOut[0][61] ), .ZN(n2554) );
  AOI22D2 U3392 ( .A1(n3400), .A2(\theRegs/completionDataOut[6][51] ), .B1(
        n3754), .B2(\theRegs/completionDataOut[7][51] ), .ZN(n2511) );
  AOI22D2 U3415 ( .A1(n3359), .A2(\theRegs/completionDataOut[4][47] ), .B1(
        n3456), .B2(\theRegs/completionDataOut[0][47] ), .ZN(n2498) );
  AOI22D2 U3485 ( .A1(n3359), .A2(\theRegs/completionDataOut[4][33] ), .B1(
        n3511), .B2(\theRegs/completionDataOut[0][33] ), .ZN(n2442) );
  AOI22D2 U3420 ( .A1(n3359), .A2(\theRegs/completionDataOut[4][46] ), .B1(
        n3493), .B2(\theRegs/completionDataOut[0][46] ), .ZN(n2494) );
  AOI22D2 U3617 ( .A1(n3374), .A2(\theRegs/completionDataOut[6][6] ), .B1(
        n4036), .B2(\theRegs/completionDataOut[7][6] ), .ZN(n2331) );
  AOI22D2 U3345 ( .A1(n3771), .A2(\theRegs/completionDataOut[4][60] ), .B1(
        n3493), .B2(\theRegs/completionDataOut[0][60] ), .ZN(n2550) );
  AOI22D2 U3378 ( .A1(n3301), .A2(\theRegs/completionDataOut[5][54] ), .B1(
        n3288), .B2(\theRegs/completionDataOut[3][54] ), .ZN(n2524) );
  AOI22D2 U3615 ( .A1(n3734), .A2(\theRegs/completionDataOut[4][7] ), .B1(
        n3511), .B2(\theRegs/completionDataOut[0][7] ), .ZN(n2338) );
  BUFFD2 U2494 ( .I(completionWriteAddr_i[2]), .Z(n3215) );
  AOI22D2 U3635 ( .A1(n3734), .A2(\theRegs/completionDataOut[4][3] ), .B1(
        n3511), .B2(\theRegs/completionDataOut[0][3] ), .ZN(n2322) );
  CKBD1 U2479 ( .I(completionWriteAddr_i[1]), .Z(n3214) );
  AOI22D2 U3450 ( .A1(n3734), .A2(\theRegs/completionDataOut[4][40] ), .B1(
        n3493), .B2(\theRegs/completionDataOut[0][40] ), .ZN(n2470) );
  INR3D1 U4125 ( .A1(n3233), .B1(n3231), .B2(n3234), .ZN(n2857) );
  BUFFD2 U3001 ( .I(n2586), .Z(n3291) );
  BUFFD2 U4193 ( .I(n2181), .Z(n3315) );
  AOI21D4 U4255 ( .A1(n3306), .A2(n2248), .B(n4027), .ZN(nextTail_o[2]) );
  BUFFD2 U4218 ( .I(n4115), .Z(n3328) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[54].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][54] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[51].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][51] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[23].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][23] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[30].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][30] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[19].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][19] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[53].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][53] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[48].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][48] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[22].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][22] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[50].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][50] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[26].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][26] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[27].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][27] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[43].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][43] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[55].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][55] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[24].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][24] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[21].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][21] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[25].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][25] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[55].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][55] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[44].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][44] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[53].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][53] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[52].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][52] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[42].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][42] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[42].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][42] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[60].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][60] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][6] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[18].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][18] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[41].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][41] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[52].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][52] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][0] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[17].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][17] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[61].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][61] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[20].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][20] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[63].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][63] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[25].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][25] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[21].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][21] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[61].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][61] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[47].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][47] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[20].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][20] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[46].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][46] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[58].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][58] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[43].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][43] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[47].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][47] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[39].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][39] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[62].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][62] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][4] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[48].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][48] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[34].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][34] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][7] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[51].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][51] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[17].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][17] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[11].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][11] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[60].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][60] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[44].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][44] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[50].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][50] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[61].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][61] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[53].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][53] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[62].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][62] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[39].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][39] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[22].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][22] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[22].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][22] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[21].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][21] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[34].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][34] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[54].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][54] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][2] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][2] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[24].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][24] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[63].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][63] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[24].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][24] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[49].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][49] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[10].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][10] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][3] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][3] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[36].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][36] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[45].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][45] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[16].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][16] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][8] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[64].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][64] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][0] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[60].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][60] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[9].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][9] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][0] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[26].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][26] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[49].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][49] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[32].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][32] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][5] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[15].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][15] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[46].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][46] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[48].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][48] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[58].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][58] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[36].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][36] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[35].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][35] ) );
  CKND2 U4835 ( .I(tail[2]), .ZN(n2265) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[22].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][22] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[33].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][33] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[35].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][35] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[64].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][64] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[38].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][38] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[23].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][23] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[37].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][37] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[59].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][59] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[31].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][31] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[33].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][33] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[52].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][52] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[40].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][40] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[28].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][28] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[10].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][10] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][1] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[32].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][32] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[37].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][37] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[31].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][31] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[27].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][27] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][5] ) );
  CKND2 U3015 ( .I(reset_i), .ZN(n2260) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[44].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][44] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[41].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][41] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[36].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][36] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[53].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][53] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[19].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][19] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[18].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][18] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[14].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][14] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][1] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[28].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][28] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][5] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[37].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][37] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[36].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][36] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[48].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][48] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][6] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[39].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][39] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][8] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[57].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][57] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[10].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][10] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[35].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][35] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][8] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][1] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[30].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][30] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[40].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][40] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[64].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][64] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[37].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][37] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[10].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][10] ) );
  INR2XD1 U3002 ( .A1(n2177), .B1(n3885), .ZN(n2179) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][6] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[14].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][14] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[28].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][28] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[53].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][53] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][2] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[37].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][37] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[29].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][29] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[15].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][15] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[49].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][49] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[45].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][45] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][4] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[9].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][9] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[26].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][26] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[12].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][12] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][2] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[29].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][29] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[52].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][52] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][1] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[34].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][34] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[35].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][35] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[27].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][27] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[64].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][64] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][5] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[44].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][44] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][6] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[45].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][45] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[30].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][30] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[16].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][16] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[12].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][12] ) );
  DFQD2 \headTailManager/tail_reg[1]  ( .D(n1401), .CP(clk_i), .Q(tail[1]) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[20].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][20] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[29].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][29] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[63].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][63] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[59].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][59] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[38].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][38] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[13].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][13] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[54].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][54] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[49].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][49] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[50].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][50] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[9].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][9] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[57].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][57] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[36].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][36] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[34].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][34] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[36].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][36] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[22].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][22] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[51].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][51] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[51].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][51] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[31].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][31] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][4] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[11].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][11] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[9].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][9] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[13].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][13] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[52].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][52] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[48].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][48] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[25].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][25] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[26].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][26] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[55].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][55] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][8] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[10].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][10] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[39].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][39] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][8] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[62].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][62] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[39].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][39] ) );
  NR3D8 U4174 ( .A1(n3246), .A2(n3240), .A3(n3241), .ZN(n2584) );
  CKND2 U2689 ( .I(n3243), .ZN(n3244) );
  ND4D8 U3611 ( .A1(n2338), .A2(n2337), .A3(n2336), .A4(n2335), .ZN(
        commitReadData_o[7]) );
  ND4D8 U3296 ( .A1(n2593), .A2(n2592), .A3(n2591), .A4(n2590), .ZN(
        commitReadData_o[69]) );
  ND4D8 U3105 ( .A1(n2310), .A2(n2309), .A3(n2308), .A4(n2307), .ZN(
        commitReadData_o[0]) );
  ND4D8 U3631 ( .A1(n2322), .A2(n2321), .A3(n2320), .A4(n2319), .ZN(
        commitReadData_o[3]) );
  NR2D2 U4178 ( .A1(n2212), .A2(n2213), .ZN(n2215) );
  CKND3 U2586 ( .I(n3225), .ZN(n3226) );
  ND4D3 U3306 ( .A1(n2578), .A2(n2577), .A3(n2576), .A4(n2575), .ZN(
        commitReadData_o[67]) );
  AOI22D2 U3522 ( .A1(n3494), .A2(\theRegs/completionDataOut[6][25] ), .B1(
        n3843), .B2(\theRegs/completionDataOut[7][25] ), .ZN(n2407) );
  AOI22D2 U3895 ( .A1(\theRegs/completionDataOut[2][13] ), .A2(n3279), .B1(
        \theRegs/completionDataOut[0][13] ), .B2(n3263), .ZN(n2806) );
  ND4D3 U3311 ( .A1(n2574), .A2(n2573), .A3(n2572), .A4(n2571), .ZN(
        commitReadData_o[66]) );
  AOI22D2 U3428 ( .A1(n3301), .A2(\theRegs/completionDataOut[5][44] ), .B1(
        n3288), .B2(\theRegs/completionDataOut[3][44] ), .ZN(n2484) );
  AOI22D2 U4019 ( .A1(\theRegs/completionDataOut[3][44] ), .A2(n3693), .B1(
        \theRegs/completionDataOut[1][44] ), .B2(n3651), .ZN(n2954) );
  AOI22D2 U3935 ( .A1(\theRegs/completionDataOut[2][5] ), .A2(n3280), .B1(
        \theRegs/completionDataOut[0][5] ), .B2(n3264), .ZN(n2838) );
  AOI22D2 U3827 ( .A1(\theRegs/completionDataOut[7][26] ), .A2(n3667), .B1(
        \theRegs/completionDataOut[6][26] ), .B2(n3716), .ZN(n2751) );
  AOI22D2 U3915 ( .A1(\theRegs/completionDataOut[2][9] ), .A2(n3280), .B1(
        \theRegs/completionDataOut[0][9] ), .B2(n3264), .ZN(n2822) );
  AOI22D2 U3880 ( .A1(\theRegs/completionDataOut[2][16] ), .A2(n3279), .B1(
        \theRegs/completionDataOut[0][16] ), .B2(n3263), .ZN(n2794) );
  AOI22D2 U3979 ( .A1(\theRegs/completionDataOut[3][37] ), .A2(n3693), .B1(
        \theRegs/completionDataOut[1][37] ), .B2(n3651), .ZN(n2982) );
  AOI22D2 U3905 ( .A1(\theRegs/completionDataOut[2][11] ), .A2(n3441), .B1(
        \theRegs/completionDataOut[0][11] ), .B2(n3410), .ZN(n2814) );
  AOI22D2 U3900 ( .A1(\theRegs/completionDataOut[2][12] ), .A2(n3441), .B1(
        \theRegs/completionDataOut[0][12] ), .B2(n3410), .ZN(n2810) );
  AOI22D2 U3143 ( .A1(\theRegs/completionDataOut[3][21] ), .A2(n3580), .B1(
        \theRegs/completionDataOut[1][21] ), .B2(n3514), .ZN(n3046) );
  AOI22D2 U3920 ( .A1(\theRegs/completionDataOut[2][8] ), .A2(n3280), .B1(
        \theRegs/completionDataOut[0][8] ), .B2(n3445), .ZN(n2826) );
  AOI22D2 U3890 ( .A1(\theRegs/completionDataOut[2][14] ), .A2(n3441), .B1(
        \theRegs/completionDataOut[0][14] ), .B2(n3410), .ZN(n2802) );
  AOI22D2 U3148 ( .A1(\theRegs/completionDataOut[3][20] ), .A2(n3580), .B1(
        \theRegs/completionDataOut[1][20] ), .B2(n3514), .ZN(n3050) );
  AOI22D2 U4102 ( .A1(\theRegs/completionDataOut[7][0] ), .A2(n3667), .B1(
        \theRegs/completionDataOut[6][0] ), .B2(n3716), .ZN(n2863) );
  AOI22D2 U3974 ( .A1(\theRegs/completionDataOut[3][36] ), .A2(n3693), .B1(
        \theRegs/completionDataOut[1][36] ), .B2(n3651), .ZN(n2986) );
  AOI22D2 U3994 ( .A1(\theRegs/completionDataOut[3][39] ), .A2(n3693), .B1(
        \theRegs/completionDataOut[1][39] ), .B2(n3651), .ZN(n2974) );
  AOI22D2 U3832 ( .A1(\theRegs/completionDataOut[7][25] ), .A2(n3667), .B1(
        \theRegs/completionDataOut[6][25] ), .B2(n3716), .ZN(n2755) );
  AOI22D2 U3964 ( .A1(\theRegs/completionDataOut[3][34] ), .A2(n3580), .B1(
        \theRegs/completionDataOut[1][34] ), .B2(n3531), .ZN(n2994) );
  AOI22D2 U3930 ( .A1(\theRegs/completionDataOut[2][6] ), .A2(n3471), .B1(
        \theRegs/completionDataOut[0][6] ), .B2(n3445), .ZN(n2834) );
  ND4D2 U3316 ( .A1(n2570), .A2(n2569), .A3(n2568), .A4(n2567), .ZN(
        commitReadData_o[65]) );
  AOI22D2 U3812 ( .A1(\theRegs/completionDataOut[7][29] ), .A2(n3667), .B1(
        \theRegs/completionDataOut[6][29] ), .B2(n3716), .ZN(n2739) );
  AOI22D2 U3774 ( .A1(\theRegs/completionDataOut[3][37] ), .A2(n3650), .B1(
        \theRegs/completionDataOut[1][37] ), .B2(n3692), .ZN(n2709) );
  AOI22D2 U3548 ( .A1(n3301), .A2(\theRegs/completionDataOut[5][20] ), .B1(
        n3287), .B2(\theRegs/completionDataOut[3][20] ), .ZN(n2388) );
  AOI22D2 U3859 ( .A1(\theRegs/completionDataOut[3][20] ), .A2(n3717), .B1(
        \theRegs/completionDataOut[1][20] ), .B2(n3671), .ZN(n2777) );
  AOI22D2 U3625 ( .A1(n3734), .A2(\theRegs/completionDataOut[4][5] ), .B1(
        n3511), .B2(\theRegs/completionDataOut[0][5] ), .ZN(n2330) );
  AOI22D2 U3885 ( .A1(\theRegs/completionDataOut[2][15] ), .A2(n3525), .B1(
        \theRegs/completionDataOut[0][15] ), .B2(n3492), .ZN(n2798) );
  AOI22D2 U3854 ( .A1(\theRegs/completionDataOut[3][21] ), .A2(n3717), .B1(
        \theRegs/completionDataOut[1][21] ), .B2(n3671), .ZN(n2773) );
  AOI22D2 U3402 ( .A1(n3405), .A2(\theRegs/completionDataOut[6][49] ), .B1(
        n3754), .B2(\theRegs/completionDataOut[7][49] ), .ZN(n2503) );
  CKBD3 U4223 ( .I(n2191), .Z(n3333) );
  AOI22D2 U3982 ( .A1(\theRegs/completionDataOut[7][64] ), .A2(n3571), .B1(
        \theRegs/completionDataOut[6][64] ), .B2(n3608), .ZN(n2599) );
  CKBD4 U4229 ( .I(n2194), .Z(n3339) );
  AOI22D2 U4105 ( .A1(\theRegs/completionDataOut[2][0] ), .A2(n3471), .B1(
        \theRegs/completionDataOut[0][0] ), .B2(n3445), .ZN(n2866) );
  AOI22D2 U3395 ( .A1(n3359), .A2(\theRegs/completionDataOut[4][51] ), .B1(
        n3493), .B2(\theRegs/completionDataOut[0][51] ), .ZN(n2514) );
  AOI22D2 U3779 ( .A1(\theRegs/completionDataOut[3][36] ), .A2(n3650), .B1(
        \theRegs/completionDataOut[1][36] ), .B2(n3692), .ZN(n2713) );
  AOI22D2 U3789 ( .A1(\theRegs/completionDataOut[3][34] ), .A2(n3717), .B1(
        \theRegs/completionDataOut[1][34] ), .B2(n3671), .ZN(n2721) );
  AOI22D2 U3453 ( .A1(n3352), .A2(\theRegs/completionDataOut[5][39] ), .B1(
        n3286), .B2(\theRegs/completionDataOut[3][39] ), .ZN(n2464) );
  AOI22D2 U3607 ( .A1(n3374), .A2(\theRegs/completionDataOut[6][8] ), .B1(
        n3843), .B2(\theRegs/completionDataOut[7][8] ), .ZN(n2339) );
  AOI22D2 U3710 ( .A1(\theRegs/completionDataOut[2][51] ), .A2(n3525), .B1(
        \theRegs/completionDataOut[0][51] ), .B2(n3492), .ZN(n2654) );
  AOI22D2 U3136 ( .A1(\theRegs/completionDataOut[7][22] ), .A2(n3368), .B1(
        \theRegs/completionDataOut[4][22] ), .B2(n3714), .ZN(n3040) );
  AOI22D2 U3128 ( .A1(\theRegs/completionDataOut[3][24] ), .A2(n3580), .B1(
        \theRegs/completionDataOut[1][24] ), .B2(n3531), .ZN(n3034) );
  AOI22D2 U3600 ( .A1(n3369), .A2(\theRegs/completionDataOut[4][10] ), .B1(
        n3511), .B2(\theRegs/completionDataOut[0][10] ), .ZN(n2350) );
  AOI22D2 U4042 ( .A1(\theRegs/completionDataOut[7][49] ), .A2(n3570), .B1(
        \theRegs/completionDataOut[4][49] ), .B2(n3532), .ZN(n2932) );
  AOI22D2 U3507 ( .A1(n3516), .A2(\theRegs/completionDataOut[6][28] ), .B1(
        n3843), .B2(\theRegs/completionDataOut[7][28] ), .ZN(n2419) );
  AOI22D2 U3839 ( .A1(\theRegs/completionDataOut[3][24] ), .A2(n3765), .B1(
        \theRegs/completionDataOut[1][24] ), .B2(n3712), .ZN(n2761) );
  AOI22D2 U3652 ( .A1(\theRegs/completionDataOut[7][48] ), .A2(n3571), .B1(
        \theRegs/completionDataOut[6][48] ), .B2(n3608), .ZN(n2663) );
  AOI22D2 U4037 ( .A1(\theRegs/completionDataOut[7][48] ), .A2(n3673), .B1(
        \theRegs/completionDataOut[4][48] ), .B2(n3629), .ZN(n2936) );
  AOI22D2 U3720 ( .A1(\theRegs/completionDataOut[2][53] ), .A2(n3525), .B1(
        \theRegs/completionDataOut[0][53] ), .B2(n3492), .ZN(n2646) );
  AOI22D2 U3670 ( .A1(\theRegs/completionDataOut[2][45] ), .A2(n3471), .B1(
        \theRegs/completionDataOut[0][45] ), .B2(n3445), .ZN(n2678) );
  AOI22D2 U3715 ( .A1(\theRegs/completionDataOut[2][52] ), .A2(n3525), .B1(
        \theRegs/completionDataOut[0][52] ), .B2(n3492), .ZN(n2650) );
  AOI22D2 U3847 ( .A1(\theRegs/completionDataOut[7][22] ), .A2(n3699), .B1(
        \theRegs/completionDataOut[6][22] ), .B2(n3744), .ZN(n2767) );
  AOI22D2 U4067 ( .A1(\theRegs/completionDataOut[7][54] ), .A2(n3673), .B1(
        \theRegs/completionDataOut[4][54] ), .B2(n3629), .ZN(n2912) );
  AOI22D2 U3829 ( .A1(\theRegs/completionDataOut[3][26] ), .A2(n3765), .B1(
        \theRegs/completionDataOut[1][26] ), .B2(n3712), .ZN(n2753) );
  AOI22D2 U3113 ( .A1(\theRegs/completionDataOut[3][27] ), .A2(n3666), .B1(
        \theRegs/completionDataOut[1][27] ), .B2(n3531), .ZN(n3022) );
  AOI22D2 U4057 ( .A1(\theRegs/completionDataOut[7][52] ), .A2(n3691), .B1(
        \theRegs/completionDataOut[4][52] ), .B2(n3649), .ZN(n2920) );
  AOI22D2 U3203 ( .A1(\theRegs/completionDataOut[3][9] ), .A2(n3666), .B1(
        \theRegs/completionDataOut[1][9] ), .B2(n3531), .ZN(n3094) );
  AOI22D2 U3817 ( .A1(\theRegs/completionDataOut[7][28] ), .A2(n3699), .B1(
        \theRegs/completionDataOut[6][28] ), .B2(n3744), .ZN(n2743) );
  AOI22D2 U3502 ( .A1(n3516), .A2(\theRegs/completionDataOut[6][29] ), .B1(
        n3843), .B2(\theRegs/completionDataOut[7][29] ), .ZN(n2423) );
  AOI22D2 U3929 ( .A1(\theRegs/completionDataOut[3][6] ), .A2(n3765), .B1(
        \theRegs/completionDataOut[1][6] ), .B2(n3712), .ZN(n2833) );
  CKBD4 U3099 ( .I(n2201), .Z(n3308) );
  AOI22D2 U3824 ( .A1(\theRegs/completionDataOut[3][27] ), .A2(n3765), .B1(
        \theRegs/completionDataOut[1][27] ), .B2(n3712), .ZN(n2749) );
  AOI22D2 U3917 ( .A1(\theRegs/completionDataOut[7][8] ), .A2(n3699), .B1(
        \theRegs/completionDataOut[6][8] ), .B2(n3744), .ZN(n2823) );
  AOI22D2 U3218 ( .A1(\theRegs/completionDataOut[3][6] ), .A2(n3666), .B1(
        \theRegs/completionDataOut[1][6] ), .B2(n3626), .ZN(n3106) );
  AOI22D2 U3463 ( .A1(n3352), .A2(\theRegs/completionDataOut[5][37] ), .B1(
        n3378), .B2(\theRegs/completionDataOut[3][37] ), .ZN(n2456) );
  AOI22D2 U3987 ( .A1(\theRegs/completionDataOut[7][38] ), .A2(n3691), .B1(
        \theRegs/completionDataOut[4][38] ), .B2(n3649), .ZN(n2976) );
  AOI22D2 U4062 ( .A1(\theRegs/completionDataOut[7][53] ), .A2(n3691), .B1(
        \theRegs/completionDataOut[4][53] ), .B2(n3649), .ZN(n2916) );
  AOI22D2 U3540 ( .A1(n3369), .A2(\theRegs/completionDataOut[4][22] ), .B1(
        n3547), .B2(\theRegs/completionDataOut[0][22] ), .ZN(n2398) );
  AOI22D2 U3206 ( .A1(\theRegs/completionDataOut[7][8] ), .A2(n3375), .B1(
        \theRegs/completionDataOut[4][8] ), .B2(n3795), .ZN(n3096) );
  AOI22D2 U3790 ( .A1(\theRegs/completionDataOut[2][34] ), .A2(n3471), .B1(
        \theRegs/completionDataOut[0][34] ), .B2(n3445), .ZN(n2722) );
  AOI22D2 U3216 ( .A1(\theRegs/completionDataOut[7][6] ), .A2(n3375), .B1(
        \theRegs/completionDataOut[4][6] ), .B2(n3795), .ZN(n3104) );
  AOI22D2 U3784 ( .A1(\theRegs/completionDataOut[3][35] ), .A2(n3650), .B1(
        \theRegs/completionDataOut[1][35] ), .B2(n3692), .ZN(n2717) );
  AOI22D2 U3618 ( .A1(n3352), .A2(\theRegs/completionDataOut[5][6] ), .B1(
        n3287), .B2(\theRegs/completionDataOut[3][6] ), .ZN(n2332) );
  AOI22D2 U3730 ( .A1(\theRegs/completionDataOut[2][55] ), .A2(n3525), .B1(
        \theRegs/completionDataOut[0][55] ), .B2(n3492), .ZN(n2638) );
  AOI22D2 U3208 ( .A1(\theRegs/completionDataOut[3][8] ), .A2(n3666), .B1(
        \theRegs/completionDataOut[1][8] ), .B2(n3626), .ZN(n3098) );
  AOI22D2 U3755 ( .A1(\theRegs/completionDataOut[2][49] ), .A2(n3544), .B1(
        \theRegs/completionDataOut[0][49] ), .B2(n3508), .ZN(n2662) );
  AOI22D2 U3934 ( .A1(\theRegs/completionDataOut[3][5] ), .A2(n3765), .B1(
        \theRegs/completionDataOut[1][5] ), .B2(n3712), .ZN(n2837) );
  AOI22D2 U3752 ( .A1(\theRegs/completionDataOut[7][49] ), .A2(n3571), .B1(
        \theRegs/completionDataOut[6][49] ), .B2(n3608), .ZN(n2659) );
  AOI22D2 U3705 ( .A1(\theRegs/completionDataOut[2][50] ), .A2(n3544), .B1(
        \theRegs/completionDataOut[0][50] ), .B2(n3508), .ZN(n2658) );
  CKBD3 U4224 ( .I(n2191), .Z(n3334) );
  CKBD3 U4230 ( .I(n2194), .Z(n3340) );
  AOI22D2 U3223 ( .A1(\theRegs/completionDataOut[3][5] ), .A2(n3698), .B1(
        \theRegs/completionDataOut[1][5] ), .B2(n3655), .ZN(n3110) );
  AOI22D2 U3196 ( .A1(\theRegs/completionDataOut[7][10] ), .A2(n3375), .B1(
        \theRegs/completionDataOut[4][10] ), .B2(n3795), .ZN(n3088) );
  INR2XD2 U4206 ( .A1(n2180), .B1(n2212), .ZN(n2181) );
  AOI22D2 U3907 ( .A1(\theRegs/completionDataOut[7][10] ), .A2(n3699), .B1(
        \theRegs/completionDataOut[6][10] ), .B2(n3744), .ZN(n2815) );
  AOI22D2 U3875 ( .A1(\theRegs/completionDataOut[2][17] ), .A2(n3544), .B1(
        \theRegs/completionDataOut[0][17] ), .B2(n3508), .ZN(n2790) );
  AOI22D2 U3528 ( .A1(n3500), .A2(\theRegs/completionDataOut[5][24] ), .B1(
        n3287), .B2(\theRegs/completionDataOut[3][24] ), .ZN(n2404) );
  CKBD4 U4158 ( .I(n2202), .Z(n3310) );
  AOI22D2 U3740 ( .A1(\theRegs/completionDataOut[2][57] ), .A2(n3544), .B1(
        \theRegs/completionDataOut[0][57] ), .B2(n3508), .ZN(n2630) );
  AOI22D2 U3914 ( .A1(\theRegs/completionDataOut[3][9] ), .A2(n3765), .B1(
        \theRegs/completionDataOut[1][9] ), .B2(n3712), .ZN(n2821) );
  AOI22D2 U3700 ( .A1(\theRegs/completionDataOut[2][39] ), .A2(n3509), .B1(
        \theRegs/completionDataOut[0][39] ), .B2(n3470), .ZN(n2702) );
  AOI22D2 U3118 ( .A1(\theRegs/completionDataOut[3][26] ), .A2(n3698), .B1(
        \theRegs/completionDataOut[1][26] ), .B2(n3655), .ZN(n3026) );
  AOI22D2 U3495 ( .A1(n3373), .A2(\theRegs/completionDataOut[4][31] ), .B1(
        n3547), .B2(\theRegs/completionDataOut[0][31] ), .ZN(n2434) );
  AOI22D2 U3608 ( .A1(n3500), .A2(\theRegs/completionDataOut[5][8] ), .B1(
        n3287), .B2(\theRegs/completionDataOut[3][8] ), .ZN(n2340) );
  AOI22D2 U3767 ( .A1(\theRegs/completionDataOut[7][38] ), .A2(n3676), .B1(
        \theRegs/completionDataOut[6][38] ), .B2(n3719), .ZN(n2703) );
  CKND2 U2599 ( .I(n3231), .ZN(n3232) );
  AOI22D2 U3655 ( .A1(\theRegs/completionDataOut[2][48] ), .A2(n3544), .B1(
        \theRegs/completionDataOut[0][48] ), .B2(n3508), .ZN(n2666) );
  AOI22D2 U3984 ( .A1(\theRegs/completionDataOut[3][64] ), .A2(n3768), .B1(
        \theRegs/completionDataOut[1][64] ), .B2(n3815), .ZN(n2601) );
  AOI22D2 U3805 ( .A1(\theRegs/completionDataOut[2][31] ), .A2(n3633), .B1(
        \theRegs/completionDataOut[0][31] ), .B2(n3595), .ZN(n2734) );
  AOI22D2 U4112 ( .A1(\theRegs/completionDataOut[7][2] ), .A2(n3838), .B1(
        \theRegs/completionDataOut[6][2] ), .B2(n3877), .ZN(n2847) );
  AOI22D2 U4117 ( .A1(\theRegs/completionDataOut[7][3] ), .A2(n3838), .B1(
        \theRegs/completionDataOut[6][3] ), .B2(n3877), .ZN(n2843) );
  AOI22D2 U3338 ( .A1(n3362), .A2(\theRegs/completionDataOut[5][61] ), .B1(
        n3545), .B2(\theRegs/completionDataOut[3][61] ), .ZN(n2552) );
  AOI22D2 U3500 ( .A1(n3373), .A2(\theRegs/completionDataOut[4][30] ), .B1(
        n3547), .B2(\theRegs/completionDataOut[0][30] ), .ZN(n2430) );
  AOI22D2 U4099 ( .A1(\theRegs/completionDataOut[3][64] ), .A2(n3816), .B1(
        \theRegs/completionDataOut[1][64] ), .B2(n3769), .ZN(n2874) );
  CKBD4 U4221 ( .I(n4005), .Z(n3331) );
  AOI22D2 U3537 ( .A1(n3516), .A2(\theRegs/completionDataOut[6][22] ), .B1(
        n3920), .B2(\theRegs/completionDataOut[7][22] ), .ZN(n2395) );
  AOI22D2 U3699 ( .A1(\theRegs/completionDataOut[3][39] ), .A2(n3768), .B1(
        \theRegs/completionDataOut[1][39] ), .B2(n3815), .ZN(n2701) );
  AOI22D2 U3919 ( .A1(\theRegs/completionDataOut[3][8] ), .A2(n3878), .B1(
        \theRegs/completionDataOut[1][8] ), .B2(n3834), .ZN(n2825) );
  AOI22D2 U3850 ( .A1(\theRegs/completionDataOut[2][22] ), .A2(n3633), .B1(
        \theRegs/completionDataOut[0][22] ), .B2(n3595), .ZN(n2770) );
  AOI22D2 U3725 ( .A1(\theRegs/completionDataOut[2][54] ), .A2(n3633), .B1(
        \theRegs/completionDataOut[0][54] ), .B2(n3595), .ZN(n2642) );
  AOI22D2 U3865 ( .A1(\theRegs/completionDataOut[2][19] ), .A2(n3705), .B1(
        \theRegs/completionDataOut[0][19] ), .B2(n3615), .ZN(n2782) );
  AOI22D2 U3717 ( .A1(\theRegs/completionDataOut[7][53] ), .A2(n3676), .B1(
        \theRegs/completionDataOut[6][53] ), .B2(n3719), .ZN(n2643) );
  AOI22D2 U3810 ( .A1(\theRegs/completionDataOut[2][30] ), .A2(n3705), .B1(
        \theRegs/completionDataOut[0][30] ), .B2(n3615), .ZN(n2738) );
  AOI22D2 U3855 ( .A1(\theRegs/completionDataOut[2][21] ), .A2(n3705), .B1(
        \theRegs/completionDataOut[0][21] ), .B2(n3615), .ZN(n2774) );
  AOI22D2 U3620 ( .A1(n3734), .A2(\theRegs/completionDataOut[4][6] ), .B1(
        n3831), .B2(\theRegs/completionDataOut[0][6] ), .ZN(n2334) );
  AOI22D2 U3972 ( .A1(\theRegs/completionDataOut[7][36] ), .A2(n3814), .B1(
        \theRegs/completionDataOut[4][36] ), .B2(n3767), .ZN(n2984) );
  AOI22D2 U3697 ( .A1(\theRegs/completionDataOut[7][39] ), .A2(n3676), .B1(
        \theRegs/completionDataOut[6][39] ), .B2(n3719), .ZN(n2699) );
  AOI22D2 U3238 ( .A1(\theRegs/completionDataOut[3][2] ), .A2(n3698), .B1(
        \theRegs/completionDataOut[1][2] ), .B2(n3655), .ZN(n3122) );
  AOI22D2 U4114 ( .A1(\theRegs/completionDataOut[3][2] ), .A2(n3878), .B1(
        \theRegs/completionDataOut[1][2] ), .B2(n3834), .ZN(n2849) );
  AOI22D2 U3775 ( .A1(\theRegs/completionDataOut[2][37] ), .A2(n3509), .B1(
        \theRegs/completionDataOut[0][37] ), .B2(n3470), .ZN(n2710) );
  AOI22D2 U3870 ( .A1(\theRegs/completionDataOut[2][18] ), .A2(n3705), .B1(
        \theRegs/completionDataOut[0][18] ), .B2(n3615), .ZN(n2786) );
  AOI22D2 U3603 ( .A1(n3500), .A2(\theRegs/completionDataOut[5][9] ), .B1(
        n3287), .B2(\theRegs/completionDataOut[3][9] ), .ZN(n2344) );
  AOI22D2 U3860 ( .A1(\theRegs/completionDataOut[2][20] ), .A2(n3705), .B1(
        \theRegs/completionDataOut[0][20] ), .B2(n3615), .ZN(n2778) );
  AOI22D2 U3375 ( .A1(n3399), .A2(\theRegs/completionDataOut[4][55] ), .B1(
        n3493), .B2(\theRegs/completionDataOut[0][55] ), .ZN(n2530) );
  AOI22D2 U3969 ( .A1(\theRegs/completionDataOut[3][35] ), .A2(n3816), .B1(
        \theRegs/completionDataOut[1][35] ), .B2(n3769), .ZN(n2990) );
  AOI22D2 U3478 ( .A1(n3362), .A2(\theRegs/completionDataOut[5][34] ), .B1(
        n3378), .B2(\theRegs/completionDataOut[3][34] ), .ZN(n2444) );
  AOI22D2 U3605 ( .A1(n3399), .A2(\theRegs/completionDataOut[4][9] ), .B1(
        n3831), .B2(\theRegs/completionDataOut[0][9] ), .ZN(n2346) );
  AOI22D2 U3939 ( .A1(\theRegs/completionDataOut[3][4] ), .A2(n3878), .B1(
        \theRegs/completionDataOut[1][4] ), .B2(n3834), .ZN(n2841) );
  AOI22D2 U3777 ( .A1(\theRegs/completionDataOut[7][36] ), .A2(n3694), .B1(
        \theRegs/completionDataOut[6][36] ), .B2(n3739), .ZN(n2711) );
  AOI22D2 U3610 ( .A1(n3399), .A2(\theRegs/completionDataOut[4][8] ), .B1(
        n3831), .B2(\theRegs/completionDataOut[0][8] ), .ZN(n2342) );
  AOI22D2 U3780 ( .A1(\theRegs/completionDataOut[2][36] ), .A2(n3509), .B1(
        \theRegs/completionDataOut[0][36] ), .B2(n3470), .ZN(n2714) );
  AOI22D2 U3228 ( .A1(\theRegs/completionDataOut[3][4] ), .A2(n3698), .B1(
        \theRegs/completionDataOut[1][4] ), .B2(n3655), .ZN(n3114) );
  AOI22D2 U3712 ( .A1(\theRegs/completionDataOut[7][52] ), .A2(n3694), .B1(
        \theRegs/completionDataOut[6][52] ), .B2(n3739), .ZN(n2647) );
  AOI22D2 U3407 ( .A1(n3405), .A2(\theRegs/completionDataOut[6][48] ), .B1(
        n3818), .B2(\theRegs/completionDataOut[7][48] ), .ZN(n2499) );
  AOI22D2 U4109 ( .A1(\theRegs/completionDataOut[3][1] ), .A2(n3878), .B1(
        \theRegs/completionDataOut[1][1] ), .B2(n3834), .ZN(n2853) );
  AOI22D2 U3468 ( .A1(n3362), .A2(\theRegs/completionDataOut[5][36] ), .B1(
        n3378), .B2(\theRegs/completionDataOut[3][36] ), .ZN(n2452) );
  AOI22D2 U3243 ( .A1(\theRegs/completionDataOut[3][1] ), .A2(n3837), .B1(
        \theRegs/completionDataOut[1][1] ), .B2(n3788), .ZN(n3126) );
  AOI22D2 U3322 ( .A1(n3405), .A2(\theRegs/completionDataOut[6][64] ), .B1(
        n3818), .B2(\theRegs/completionDataOut[7][64] ), .ZN(n2563) );
  AOI22D2 U3387 ( .A1(n3405), .A2(\theRegs/completionDataOut[6][52] ), .B1(
        n3818), .B2(\theRegs/completionDataOut[7][52] ), .ZN(n2515) );
  OAI21D4 U4168 ( .A1(tailReset), .A2(n2269), .B(n2260), .ZN(n2264) );
  AOI22D2 U3373 ( .A1(n3641), .A2(\theRegs/completionDataOut[5][55] ), .B1(
        n3545), .B2(\theRegs/completionDataOut[3][55] ), .ZN(n2528) );
  AOI22D2 U3380 ( .A1(n3579), .A2(\theRegs/completionDataOut[4][54] ), .B1(
        n3493), .B2(\theRegs/completionDataOut[0][54] ), .ZN(n2526) );
  AOI22D2 U3385 ( .A1(n3579), .A2(\theRegs/completionDataOut[4][53] ), .B1(
        n3515), .B2(\theRegs/completionDataOut[0][53] ), .ZN(n2522) );
  AOI22D2 U3323 ( .A1(n3362), .A2(\theRegs/completionDataOut[5][64] ), .B1(
        n3378), .B2(\theRegs/completionDataOut[3][64] ), .ZN(n2564) );
  AOI22D2 U3597 ( .A1(n3374), .A2(\theRegs/completionDataOut[6][10] ), .B1(
        n3920), .B2(\theRegs/completionDataOut[7][10] ), .ZN(n2347) );
  AOI22D2 U3543 ( .A1(n3641), .A2(\theRegs/completionDataOut[5][21] ), .B1(
        n3350), .B2(\theRegs/completionDataOut[3][21] ), .ZN(n2392) );
  AOI22D2 U3382 ( .A1(n3405), .A2(\theRegs/completionDataOut[6][53] ), .B1(
        n3818), .B2(\theRegs/completionDataOut[7][53] ), .ZN(n2519) );
  AOI22D2 U3513 ( .A1(n3641), .A2(\theRegs/completionDataOut[5][27] ), .B1(
        n3350), .B2(\theRegs/completionDataOut[3][27] ), .ZN(n2416) );
  INR2XD2 U3051 ( .A1(n2213), .B1(n2212), .ZN(n2214) );
  AOI22D2 U3405 ( .A1(n3579), .A2(\theRegs/completionDataOut[4][49] ), .B1(
        n3515), .B2(\theRegs/completionDataOut[0][49] ), .ZN(n2506) );
  AOI22D2 U3390 ( .A1(n3579), .A2(\theRegs/completionDataOut[4][52] ), .B1(
        n3515), .B2(\theRegs/completionDataOut[0][52] ), .ZN(n2518) );
  AOI22D2 U3518 ( .A1(n3682), .A2(\theRegs/completionDataOut[5][26] ), .B1(
        n3350), .B2(\theRegs/completionDataOut[3][26] ), .ZN(n2412) );
  AOI22D2 U3365 ( .A1(n3579), .A2(\theRegs/completionDataOut[4][57] ), .B1(
        n3515), .B2(\theRegs/completionDataOut[0][57] ), .ZN(n2538) );
  AOI22D2 U3410 ( .A1(n3579), .A2(\theRegs/completionDataOut[4][48] ), .B1(
        n3534), .B2(\theRegs/completionDataOut[0][48] ), .ZN(n2502) );
  AOI22D2 U3623 ( .A1(n3362), .A2(\theRegs/completionDataOut[5][5] ), .B1(
        n3350), .B2(\theRegs/completionDataOut[3][5] ), .ZN(n2328) );
  AOI22D2 U3638 ( .A1(n3366), .A2(\theRegs/completionDataOut[5][2] ), .B1(
        n3378), .B2(\theRegs/completionDataOut[3][2] ), .ZN(n2316) );
  AOI22D2 U3470 ( .A1(n3734), .A2(\theRegs/completionDataOut[4][36] ), .B1(
        n3534), .B2(\theRegs/completionDataOut[0][36] ), .ZN(n2454) );
  INR2XD2 U3098 ( .A1(n2228), .B1(n2229), .ZN(n2231) );
  AOI22D2 U3465 ( .A1(n3597), .A2(\theRegs/completionDataOut[4][37] ), .B1(
        n3534), .B2(\theRegs/completionDataOut[0][37] ), .ZN(n2458) );
  INR2XD1 U2805 ( .A1(n2183), .B1(n2216), .ZN(n2184) );
  AOI22D2 U3628 ( .A1(n3366), .A2(\theRegs/completionDataOut[5][4] ), .B1(
        n3386), .B2(\theRegs/completionDataOut[3][4] ), .ZN(n2324) );
  NR2D2 U4164 ( .A1(n2216), .A2(n2183), .ZN(n2185) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[57].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][57] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[17].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][17] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[56].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][56] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[21].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[21].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][21] ) );
  CKND2 U4834 ( .I(tail[1]), .ZN(n2262) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[13].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][13] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[16].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][16] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[27].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][27] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[50].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][50] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[15].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][15] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[14].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][14] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[34].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][34] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[56].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][56] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[23].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][23] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[31].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][31] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[24].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][24] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[34].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][34] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[51].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][51] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[11].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][11] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][3] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[41].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][41] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[42].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][42] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][4] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[27].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][27] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[58].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][58] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][7] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[12].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][12] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[24].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][24] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[9].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][9] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[19].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][19] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[10].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][10] ) );
  INR2XD1 U2867 ( .A1(n3372), .B1(n2236), .ZN(n2197) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][1] ) );
  CKBD3 U4220 ( .I(n2187), .Z(n3330) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[56].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][56] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][2] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[11].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][11] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[16].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][16] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[33].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][33] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[44].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][44] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[57].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][57] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[45].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][45] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[50].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][50] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[41].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][41] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[29].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][29] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[23].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][23] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[28].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][28] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[30].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][30] ) );
  IND2D1 U4824 ( .A1(n2247), .B1(n2243), .ZN(n2233) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[9].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][9] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[20].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][20] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[64].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][64] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[51].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][51] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[15].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][15] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[33].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][33] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[32].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][32] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[41].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][41] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[30].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][30] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[40].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][40] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[43].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][43] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[43].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][43] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[35].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][35] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[25].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][25] ) );
  AOI22D4 U3294 ( .A1(n3683), .A2(\theRegs/managementDataOut[1][0] ), .B1(
        n3831), .B2(\theRegs/managementDataOut[0][0] ), .ZN(n2273) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[52].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][52] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][3] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[55].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][55] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[43].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][43] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[13].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][13] ) );
  AOI22D4 U3295 ( .A1(n3366), .A2(\theRegs/managementDataOut[5][0] ), .B1(
        n3597), .B2(\theRegs/managementDataOut[4][0] ), .ZN(n2274) );
  AOI22D4 U3284 ( .A1(n3855), .A2(\theRegs/managementDataOut[1][2] ), .B1(
        n3831), .B2(\theRegs/managementDataOut[0][2] ), .ZN(n2281) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[42].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][42] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[58].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][58] ) );
  NR3D4 U4180 ( .A1(n3242), .A2(n3240), .A3(n3245), .ZN(n2589) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][7] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[32].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][32] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[41].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][41] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[14].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][14] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[40].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][40] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[18].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][18] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[62].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][62] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[23].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][23] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[59].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][59] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[43].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][43] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[40].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][40] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[58].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][58] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[46].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][46] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[47].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][47] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[56].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][56] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[60].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][60] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][7] ) );
  OAI221D4 U2288 ( .A1(n3240), .A2(n2207), .B1(n3242), .B2(n3283), .C(n2204), 
        .ZN(n2206) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[32].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][32] ) );
  CKBD3 U2475 ( .I(completionWriteAddr_i[0]), .Z(n3212) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[45].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][45] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[45].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][45] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[12].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][12] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[57].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][57] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[59].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][59] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[58].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][58] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[31].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][31] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[60].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][60] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][3] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[46].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][46] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[33].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][33] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[48].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][48] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[33].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][33] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[51].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][51] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[46].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][46] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[22].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][22] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[54].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][54] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[33].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][33] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[17].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][17] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[42].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][42] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[62].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][62] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[50].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][50] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[53].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][53] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[17].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[17].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][17] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[59].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][59] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[22].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][22] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[10].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[10].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][10] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[47].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][47] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[46].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][46] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[63].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][63] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[23].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][23] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[56].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][56] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[55].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][55] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[40].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][40] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[54].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][54] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[29].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][29] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[64].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][64] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[23].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][23] ) );
  AOI22D4 U3280 ( .A1(n3366), .A2(\theRegs/managementDataOut[5][3] ), .B1(
        n3597), .B2(\theRegs/managementDataOut[4][3] ), .ZN(n2286) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[49].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][49] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[44].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][44] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[61].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][61] ) );
  AOI22D4 U3289 ( .A1(n3855), .A2(\theRegs/managementDataOut[1][1] ), .B1(
        n3831), .B2(\theRegs/managementDataOut[0][1] ), .ZN(n2277) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[54].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[54].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][54] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[49].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][49] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][4] ) );
  AOI22D4 U3279 ( .A1(n3855), .A2(\theRegs/managementDataOut[1][3] ), .B1(
        n3750), .B2(\theRegs/managementDataOut[0][3] ), .ZN(n2285) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[24].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][24] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[25].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][25] ) );
  AOI22D4 U3259 ( .A1(n3855), .A2(\theRegs/managementDataOut[1][7] ), .B1(
        n3750), .B2(\theRegs/managementDataOut[0][7] ), .ZN(n2301) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[30].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][30] ) );
  AOI22D4 U3269 ( .A1(n3967), .A2(\theRegs/managementDataOut[1][5] ), .B1(
        n3750), .B2(\theRegs/managementDataOut[0][5] ), .ZN(n2293) );
  DFQD2 \headTailManager/head_reg[1]  ( .D(n1405), .CP(clk_i), .Q(head[1]) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[38].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][38] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[32].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][32] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[26].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][26] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[58].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][58] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[63].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][63] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[59].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][59] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[42].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][42] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[47].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][47] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[38].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][38] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[43].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][43] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[19].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[19].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][19] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[15].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][15] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][5] ) );
  AOI22D4 U3304 ( .A1(n3429), .A2(\theRegs/completionDataOut[1][68] ), .B1(
        n3668), .B2(\theRegs/completionDataOut[0][68] ), .ZN(n2581) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[27].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][27] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[29].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][29] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[56].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[56].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][56] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[38].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][38] ) );
  AOI22D4 U3274 ( .A1(n3967), .A2(\theRegs/managementDataOut[1][4] ), .B1(
        n3933), .B2(\theRegs/managementDataOut[0][4] ), .ZN(n2289) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[51].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[51].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][51] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[18].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[18].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][18] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[50].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][50] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[42].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][42] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][1] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[16].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][16] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][3] ) );
  AOI22D4 U3290 ( .A1(n3517), .A2(\theRegs/managementDataOut[5][1] ), .B1(
        n3597), .B2(\theRegs/managementDataOut[4][1] ), .ZN(n2278) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[37].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][37] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[52].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][52] ) );
  DFQD2 \theRegs/eachCompletionReg[1].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[1].completionReg/eachEnDff[61].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[1][61] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[32].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][32] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[41].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][41] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[28].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][28] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[31].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][31] ) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][7] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[63].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][63] ) );
  DFQD2 \theRegs/eachCompletionReg[5].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[5].completionReg/eachEnDff[38].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[5][38] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[39].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][39] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][5] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[28].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][28] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[34].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][34] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[25].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][25] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[23].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[23].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][23] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[42].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[42].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][42] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][0] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[63].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][63] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][0] ) );
  AOI22D4 U3260 ( .A1(n3517), .A2(\theRegs/managementDataOut[5][7] ), .B1(
        n3597), .B2(\theRegs/managementDataOut[4][7] ), .ZN(n2302) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[48].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][48] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[40].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][40] ) );
  AOI22D4 U3305 ( .A1(n3517), .A2(\theRegs/completionDataOut[5][68] ), .B1(
        n3560), .B2(\theRegs/completionDataOut[4][68] ), .ZN(n2582) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[13].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][13] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[38].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[38].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][38] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][2] ) );
  BUFFD2 U2628 ( .I(decodeReadAddr1_i[1]), .Z(n3233) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[33].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[33].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][33] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[43].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[43].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][43] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[45].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][45] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[50].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[50].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][50] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[14].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][14] ) );
  AOI22D2 U3285 ( .A1(n3646), .A2(\theRegs/managementDataOut[5][2] ), .B1(
        n3560), .B2(\theRegs/managementDataOut[4][2] ), .ZN(n2282) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[58].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[58].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][58] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][7] ) );
  AOI22D4 U3255 ( .A1(\theRegs/managementDataOut[5][8] ), .A2(n3646), .B1(
        \theRegs/managementDataOut[4][8] ), .B2(n3560), .ZN(n2306) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[60].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][60] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[29].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][29] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[40].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[40].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][40] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[12].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][12] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[45].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[45].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][45] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[59].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][59] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[30].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][30] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[11].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[11].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][11] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[32].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[32].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][32] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[41].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[41].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][41] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[53].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][53] ) );
  AOI22D2 U3264 ( .A1(n3967), .A2(\theRegs/managementDataOut[1][6] ), .B1(
        n3933), .B2(\theRegs/managementDataOut[0][6] ), .ZN(n2297) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[62].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][62] ) );
  AOI22D4 U3275 ( .A1(n3646), .A2(\theRegs/managementDataOut[5][4] ), .B1(
        n3560), .B2(\theRegs/managementDataOut[4][4] ), .ZN(n2290) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[47].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][47] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[46].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][46] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[57].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][57] ) );
  DFQD4 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[16].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[16].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][16] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[31].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][31] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[62].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][62] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][7] ) );
  DFQD2 \theRegs/eachCompletionReg[2].completionReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[2].completionReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[2][3] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[60].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][60] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[37].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][37] ) );
  DFQD4 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[14].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[14].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][14] ) );
  DFQD4 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[12].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][12] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[25].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][25] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[47].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][47] ) );
  NR2XD3 U2286 ( .A1(n2270), .A2(n2269), .ZN(n2268) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[62].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[62].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][62] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[55].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][55] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[61].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][61] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[35].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][35] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[63].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[63].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][63] ) );
  DFQD4 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[15].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[15].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][15] ) );
  DFQD4 \headTailManager/tail_reg[0]  ( .D(n1402), .CP(clk_i), .Q(tail[0]) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[59].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[59].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][59] ) );
  AO22D1 U2570 ( .A1(n3194), .A2(n3985), .B1(n3807), .B2(
        \theRegs/completionDataOut[6][53] ), .Z(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[53].enDff/theFlop/N3 ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[61].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][61] ) );
  DFQD4 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[13].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[13].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][13] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[44].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][44] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[60].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[60].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][60] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[46].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[46].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][46] ) );
  DFQD4 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[12].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[12].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][12] ) );
  ND4D8 U3471 ( .A1(n2450), .A2(n2449), .A3(n2448), .A4(n2447), .ZN(
        commitReadData_o[35]) );
  ND4D8 U3636 ( .A1(n2318), .A2(n2317), .A3(n2316), .A4(n2315), .ZN(
        commitReadData_o[2]) );
  DFQD4 \headTailManager/tailReset_reg  ( .D(n1403), .CP(clk_i), .Q(tailReset)
         );
  AOI22D2 U3940 ( .A1(\theRegs/completionDataOut[2][4] ), .A2(n3509), .B1(
        \theRegs/completionDataOut[0][4] ), .B2(n3470), .ZN(n2842) );
  AOI22D2 U4110 ( .A1(\theRegs/completionDataOut[2][1] ), .A2(n3509), .B1(
        \theRegs/completionDataOut[0][1] ), .B2(n3470), .ZN(n2854) );
  AOI22D2 U4115 ( .A1(\theRegs/completionDataOut[2][2] ), .A2(n3599), .B1(
        \theRegs/completionDataOut[0][2] ), .B2(n3556), .ZN(n2850) );
  AOI22D2 U3423 ( .A1(n3682), .A2(\theRegs/completionDataOut[5][45] ), .B1(
        n3545), .B2(\theRegs/completionDataOut[3][45] ), .ZN(n2488) );
  CKND3 U2458 ( .I(completionWriteEn_i), .ZN(n3211) );
  AOI22D2 U3438 ( .A1(n3718), .A2(\theRegs/completionDataOut[5][42] ), .B1(
        n3545), .B2(\theRegs/completionDataOut[3][42] ), .ZN(n2476) );
  AOI22D2 U4052 ( .A1(\theRegs/completionDataOut[7][51] ), .A2(n3814), .B1(
        \theRegs/completionDataOut[4][51] ), .B2(n3767), .ZN(n2924) );
  AOI22D2 U3327 ( .A1(n3449), .A2(\theRegs/completionDataOut[6][63] ), .B1(
        n3841), .B2(\theRegs/completionDataOut[7][63] ), .ZN(n2559) );
  AOI22D2 U3433 ( .A1(n3718), .A2(\theRegs/completionDataOut[5][43] ), .B1(
        n3545), .B2(\theRegs/completionDataOut[3][43] ), .ZN(n2480) );
  AOI22D2 U3613 ( .A1(n3682), .A2(\theRegs/completionDataOut[5][7] ), .B1(
        n3386), .B2(\theRegs/completionDataOut[3][7] ), .ZN(n2336) );
  AOI22D2 U3201 ( .A1(\theRegs/completionDataOut[7][9] ), .A2(n3375), .B1(
        \theRegs/completionDataOut[4][9] ), .B2(n3795), .ZN(n3092) );
  AOI22D2 U3328 ( .A1(n3830), .A2(\theRegs/completionDataOut[5][63] ), .B1(
        n3402), .B2(\theRegs/completionDataOut[3][63] ), .ZN(n2560) );
  AOI22D2 U3332 ( .A1(n3462), .A2(\theRegs/completionDataOut[6][62] ), .B1(
        n3841), .B2(\theRegs/completionDataOut[7][62] ), .ZN(n2555) );
  AOI22D2 U3343 ( .A1(n3830), .A2(\theRegs/completionDataOut[5][60] ), .B1(
        n3601), .B2(\theRegs/completionDataOut[3][60] ), .ZN(n2548) );
  AOI22D2 U3947 ( .A1(\theRegs/completionDataOut[7][31] ), .A2(n3375), .B1(
        \theRegs/completionDataOut[4][31] ), .B2(n3795), .ZN(n3004) );
  AOI22D2 U3680 ( .A1(\theRegs/completionDataOut[2][43] ), .A2(n3599), .B1(
        \theRegs/completionDataOut[0][43] ), .B2(n3556), .ZN(n2686) );
  AOI22D2 U3221 ( .A1(\theRegs/completionDataOut[7][5] ), .A2(n3404), .B1(
        \theRegs/completionDataOut[4][5] ), .B2(n3880), .ZN(n3108) );
  AOI22D2 U3647 ( .A1(\theRegs/completionDataOut[7][63] ), .A2(n3694), .B1(
        \theRegs/completionDataOut[6][63] ), .B2(n3739), .ZN(n2603) );
  AOI22D2 U3400 ( .A1(n3644), .A2(\theRegs/completionDataOut[4][50] ), .B1(
        n3668), .B2(\theRegs/completionDataOut[0][50] ), .ZN(n2510) );
  AOI22D2 U3685 ( .A1(\theRegs/completionDataOut[2][42] ), .A2(n3599), .B1(
        \theRegs/completionDataOut[0][42] ), .B2(n3556), .ZN(n2690) );
  AOI22D2 U3942 ( .A1(\theRegs/completionDataOut[7][30] ), .A2(n3404), .B1(
        \theRegs/completionDataOut[4][30] ), .B2(n3880), .ZN(n3008) );
  AOI22D2 U3333 ( .A1(n3830), .A2(\theRegs/completionDataOut[5][62] ), .B1(
        n3402), .B2(\theRegs/completionDataOut[3][62] ), .ZN(n2556) );
  AOI22D2 U3418 ( .A1(n3682), .A2(\theRegs/completionDataOut[5][46] ), .B1(
        n3601), .B2(\theRegs/completionDataOut[3][46] ), .ZN(n2492) );
  AOI22D2 U3443 ( .A1(n3830), .A2(\theRegs/completionDataOut[5][41] ), .B1(
        n3402), .B2(\theRegs/completionDataOut[3][41] ), .ZN(n2472) );
  AOI22D2 U3533 ( .A1(n3682), .A2(\theRegs/completionDataOut[5][23] ), .B1(
        n3390), .B2(\theRegs/completionDataOut[3][23] ), .ZN(n2400) );
  AOI22D2 U3337 ( .A1(n3462), .A2(\theRegs/completionDataOut[6][61] ), .B1(
        n3909), .B2(\theRegs/completionDataOut[7][61] ), .ZN(n2551) );
  AOI22D2 U3785 ( .A1(\theRegs/completionDataOut[2][35] ), .A2(n3620), .B1(
        \theRegs/completionDataOut[0][35] ), .B2(n3583), .ZN(n2718) );
  AOI22D2 U4122 ( .A1(\theRegs/completionDataOut[7][60] ), .A2(n3817), .B1(
        \theRegs/completionDataOut[6][60] ), .B2(n3861), .ZN(n2615) );
  AOI22D2 U3578 ( .A1(n3707), .A2(\theRegs/completionDataOut[5][14] ), .B1(
        n3390), .B2(\theRegs/completionDataOut[3][14] ), .ZN(n2364) );
  AOI22D2 U3757 ( .A1(\theRegs/completionDataOut[7][61] ), .A2(n3817), .B1(
        \theRegs/completionDataOut[6][61] ), .B2(n3861), .ZN(n2611) );
  AOI22D2 U3408 ( .A1(n3707), .A2(\theRegs/completionDataOut[5][48] ), .B1(
        n3601), .B2(\theRegs/completionDataOut[3][48] ), .ZN(n2500) );
  AOI22D2 U3650 ( .A1(\theRegs/completionDataOut[2][63] ), .A2(n3620), .B1(
        \theRegs/completionDataOut[0][63] ), .B2(n3583), .ZN(n2606) );
  AOI22D2 U3782 ( .A1(\theRegs/completionDataOut[7][35] ), .A2(n3817), .B1(
        \theRegs/completionDataOut[6][35] ), .B2(n3861), .ZN(n2715) );
  AOI22D2 U3762 ( .A1(\theRegs/completionDataOut[7][62] ), .A2(n3817), .B1(
        \theRegs/completionDataOut[6][62] ), .B2(n3861), .ZN(n2607) );
  AOI22D2 U3985 ( .A1(\theRegs/completionDataOut[2][64] ), .A2(n3620), .B1(
        \theRegs/completionDataOut[0][64] ), .B2(n3583), .ZN(n2602) );
  AOI22D2 U3665 ( .A1(\theRegs/completionDataOut[2][46] ), .A2(n3620), .B1(
        \theRegs/completionDataOut[0][46] ), .B2(n3583), .ZN(n2674) );
  AOI22D2 U3760 ( .A1(\theRegs/completionDataOut[2][61] ), .A2(n3720), .B1(
        \theRegs/completionDataOut[0][61] ), .B2(n3672), .ZN(n2614) );
  AOI22D2 U3413 ( .A1(n3707), .A2(\theRegs/completionDataOut[5][47] ), .B1(
        n3601), .B2(\theRegs/completionDataOut[3][47] ), .ZN(n2496) );
  AOI22D2 U4072 ( .A1(\theRegs/completionDataOut[7][55] ), .A2(n3814), .B1(
        \theRegs/completionDataOut[4][55] ), .B2(n3767), .ZN(n2908) );
  AOI22D2 U3795 ( .A1(\theRegs/completionDataOut[2][33] ), .A2(n3772), .B1(
        \theRegs/completionDataOut[0][33] ), .B2(n3670), .ZN(n2726) );
  AOI22D2 U3363 ( .A1(n3707), .A2(\theRegs/completionDataOut[5][57] ), .B1(
        n3601), .B2(\theRegs/completionDataOut[3][57] ), .ZN(n2536) );
  CKBD4 U2799 ( .I(n3133), .Z(n3253) );
  AOI22D2 U3398 ( .A1(n3707), .A2(\theRegs/completionDataOut[5][50] ), .B1(
        n3654), .B2(\theRegs/completionDataOut[3][50] ), .ZN(n2508) );
  AOI22D2 U3660 ( .A1(\theRegs/completionDataOut[2][47] ), .A2(n3772), .B1(
        \theRegs/completionDataOut[0][47] ), .B2(n3670), .ZN(n2670) );
  AOI22D2 U4107 ( .A1(\theRegs/completionDataOut[7][1] ), .A2(n3838), .B1(
        \theRegs/completionDataOut[6][1] ), .B2(n3877), .ZN(n2851) );
  CKBD4 U2802 ( .I(n3132), .Z(n3255) );
  AOI22D2 U3690 ( .A1(\theRegs/completionDataOut[2][41] ), .A2(n3720), .B1(
        \theRegs/completionDataOut[0][41] ), .B2(n3672), .ZN(n2694) );
  AOI22D2 U3745 ( .A1(\theRegs/completionDataOut[2][58] ), .A2(n3772), .B1(
        \theRegs/completionDataOut[0][58] ), .B2(n3672), .ZN(n2626) );
  AOI22D2 U3800 ( .A1(\theRegs/completionDataOut[2][32] ), .A2(n3720), .B1(
        \theRegs/completionDataOut[0][32] ), .B2(n3670), .ZN(n2730) );
  AOI22D2 U3750 ( .A1(\theRegs/completionDataOut[2][59] ), .A2(n3720), .B1(
        \theRegs/completionDataOut[0][59] ), .B2(n3672), .ZN(n2622) );
  AOI22D2 U3448 ( .A1(n3830), .A2(\theRegs/completionDataOut[5][40] ), .B1(
        n3402), .B2(\theRegs/completionDataOut[3][40] ), .ZN(n2468) );
  AOI22D2 U3765 ( .A1(\theRegs/completionDataOut[2][62] ), .A2(n3746), .B1(
        \theRegs/completionDataOut[0][62] ), .B2(n3697), .ZN(n2610) );
  AOI22D2 U4127 ( .A1(\theRegs/completionDataOut[2][60] ), .A2(n3746), .B1(
        \theRegs/completionDataOut[0][60] ), .B2(n3697), .ZN(n2618) );
  AOI22D2 U3830 ( .A1(\theRegs/completionDataOut[2][26] ), .A2(n3800), .B1(
        \theRegs/completionDataOut[0][26] ), .B2(n3745), .ZN(n2754) );
  AOI22D2 U3840 ( .A1(\theRegs/completionDataOut[2][24] ), .A2(n3800), .B1(
        \theRegs/completionDataOut[0][24] ), .B2(n3745), .ZN(n2762) );
  AOI22D2 U3695 ( .A1(\theRegs/completionDataOut[2][40] ), .A2(n3746), .B1(
        \theRegs/completionDataOut[0][40] ), .B2(n3697), .ZN(n2698) );
  AOI22D2 U3825 ( .A1(\theRegs/completionDataOut[2][27] ), .A2(n3930), .B1(
        \theRegs/completionDataOut[0][27] ), .B2(n3879), .ZN(n2750) );
  AOI22D2 U3342 ( .A1(n3462), .A2(\theRegs/completionDataOut[6][60] ), .B1(
        n3909), .B2(\theRegs/completionDataOut[7][60] ), .ZN(n2547) );
  AOI22D2 U3835 ( .A1(\theRegs/completionDataOut[2][25] ), .A2(n3930), .B1(
        \theRegs/completionDataOut[0][25] ), .B2(n3879), .ZN(n2758) );
  AOI22D2 U3977 ( .A1(\theRegs/completionDataOut[7][37] ), .A2(n3814), .B1(
        \theRegs/completionDataOut[4][37] ), .B2(n3767), .ZN(n2980) );
  AOI22D2 U3508 ( .A1(n3707), .A2(\theRegs/completionDataOut[5][28] ), .B1(
        n3390), .B2(\theRegs/completionDataOut[3][28] ), .ZN(n2420) );
  AOI22D2 U3553 ( .A1(n3820), .A2(\theRegs/completionDataOut[5][19] ), .B1(
        n3390), .B2(\theRegs/completionDataOut[3][19] ), .ZN(n2384) );
  BUFFD6 U2863 ( .I(n2860), .Z(n3266) );
  AOI22D2 U3348 ( .A1(n3830), .A2(\theRegs/completionDataOut[5][59] ), .B1(
        n3654), .B2(\theRegs/completionDataOut[3][59] ), .ZN(n2544) );
  AOI22D2 U3568 ( .A1(n3820), .A2(\theRegs/completionDataOut[5][16] ), .B1(
        n3390), .B2(\theRegs/completionDataOut[3][16] ), .ZN(n2372) );
  AOI22D2 U3815 ( .A1(\theRegs/completionDataOut[2][29] ), .A2(n3930), .B1(
        \theRegs/completionDataOut[0][29] ), .B2(n3879), .ZN(n2742) );
  AOI22D2 U3820 ( .A1(\theRegs/completionDataOut[2][28] ), .A2(n3930), .B1(
        \theRegs/completionDataOut[0][28] ), .B2(n3879), .ZN(n2746) );
  BUFFD6 U2806 ( .I(n3975), .Z(n3258) );
  AOI22D2 U3523 ( .A1(n3856), .A2(\theRegs/completionDataOut[5][25] ), .B1(
        n3390), .B2(\theRegs/completionDataOut[3][25] ), .ZN(n2408) );
  CKBD4 U2800 ( .I(n3133), .Z(n3254) );
  CKBD4 U2803 ( .I(n3132), .Z(n3256) );
  AOI22D2 U3845 ( .A1(\theRegs/completionDataOut[2][23] ), .A2(n3930), .B1(
        \theRegs/completionDataOut[0][23] ), .B2(n3879), .ZN(n2766) );
  AOI22D2 U3573 ( .A1(n3856), .A2(\theRegs/completionDataOut[5][15] ), .B1(
        n3431), .B2(\theRegs/completionDataOut[3][15] ), .ZN(n2368) );
  AOI22D2 U3488 ( .A1(n3856), .A2(\theRegs/completionDataOut[5][32] ), .B1(
        n3431), .B2(\theRegs/completionDataOut[3][32] ), .ZN(n2436) );
  AOI22D2 U3598 ( .A1(n3856), .A2(\theRegs/completionDataOut[5][10] ), .B1(
        n3431), .B2(\theRegs/completionDataOut[3][10] ), .ZN(n2348) );
  AOI22D2 U3503 ( .A1(n3856), .A2(\theRegs/completionDataOut[5][29] ), .B1(
        n3431), .B2(\theRegs/completionDataOut[3][29] ), .ZN(n2424) );
  AOI22D2 U3558 ( .A1(n3908), .A2(\theRegs/completionDataOut[5][18] ), .B1(
        n3431), .B2(\theRegs/completionDataOut[3][18] ), .ZN(n2380) );
  AOI22D2 U3393 ( .A1(n3908), .A2(\theRegs/completionDataOut[5][51] ), .B1(
        n3654), .B2(\theRegs/completionDataOut[3][51] ), .ZN(n2512) );
  AOI22D2 U3388 ( .A1(n3908), .A2(\theRegs/completionDataOut[5][52] ), .B1(
        n3654), .B2(\theRegs/completionDataOut[3][52] ), .ZN(n2516) );
  AOI22D2 U3633 ( .A1(n3505), .A2(\theRegs/completionDataOut[5][3] ), .B1(
        n3481), .B2(\theRegs/completionDataOut[3][3] ), .ZN(n2320) );
  AOI22D2 U3480 ( .A1(n3466), .A2(\theRegs/completionDataOut[4][34] ), .B1(
        n3933), .B2(\theRegs/completionDataOut[0][34] ), .ZN(n2446) );
  AOI22D2 U3483 ( .A1(n3908), .A2(\theRegs/completionDataOut[5][33] ), .B1(
        n3778), .B2(\theRegs/completionDataOut[3][33] ), .ZN(n2440) );
  AOI22D2 U3498 ( .A1(n3951), .A2(\theRegs/completionDataOut[5][30] ), .B1(
        n3530), .B2(\theRegs/completionDataOut[3][30] ), .ZN(n2428) );
  AOI22D2 U3563 ( .A1(n3951), .A2(\theRegs/completionDataOut[5][17] ), .B1(
        n3530), .B2(\theRegs/completionDataOut[3][17] ), .ZN(n2376) );
  AOI22D2 U3583 ( .A1(n3951), .A2(\theRegs/completionDataOut[5][13] ), .B1(
        n3530), .B2(\theRegs/completionDataOut[3][13] ), .ZN(n2360) );
  AOI22D2 U3538 ( .A1(n3951), .A2(\theRegs/completionDataOut[5][22] ), .B1(
        n3530), .B2(\theRegs/completionDataOut[3][22] ), .ZN(n2396) );
  AOI22D2 U3493 ( .A1(n3951), .A2(\theRegs/completionDataOut[5][31] ), .B1(
        n3530), .B2(\theRegs/completionDataOut[3][31] ), .ZN(n2432) );
  AOI22D2 U3383 ( .A1(n4004), .A2(\theRegs/completionDataOut[5][53] ), .B1(
        n3778), .B2(\theRegs/completionDataOut[3][53] ), .ZN(n2520) );
  AOI22D2 U3588 ( .A1(n4004), .A2(\theRegs/completionDataOut[5][12] ), .B1(
        n3591), .B2(\theRegs/completionDataOut[3][12] ), .ZN(n2356) );
  AOI22D2 U3593 ( .A1(n4004), .A2(\theRegs/completionDataOut[5][11] ), .B1(
        n3591), .B2(\theRegs/completionDataOut[3][11] ), .ZN(n2352) );
  AOI22D2 U3353 ( .A1(n4004), .A2(\theRegs/completionDataOut[5][58] ), .B1(
        n3778), .B2(\theRegs/completionDataOut[3][58] ), .ZN(n2540) );
  AOI22D2 U3430 ( .A1(n3644), .A2(\theRegs/completionDataOut[4][44] ), .B1(
        n3668), .B2(\theRegs/completionDataOut[0][44] ), .ZN(n2486) );
  AOI22D2 U3107 ( .A1(n3505), .A2(\theRegs/completionDataOut[5][0] ), .B1(
        n3402), .B2(\theRegs/completionDataOut[3][0] ), .ZN(n2308) );
  AOI22D2 U3425 ( .A1(n3644), .A2(\theRegs/completionDataOut[4][45] ), .B1(
        n3801), .B2(\theRegs/completionDataOut[0][45] ), .ZN(n2490) );
  AOI22D2 U3455 ( .A1(n3466), .A2(\theRegs/completionDataOut[4][39] ), .B1(
        n3801), .B2(\theRegs/completionDataOut[0][39] ), .ZN(n2466) );
  CKBD4 U3063 ( .I(\add_x_7/n1 ), .Z(n3302) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[53].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[53].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][53] ) );
  AOI22D2 U3460 ( .A1(n3466), .A2(\theRegs/completionDataOut[4][38] ), .B1(
        n3801), .B2(\theRegs/completionDataOut[0][38] ), .ZN(n2462) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][8] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[20].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[20].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][20] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[52].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[52].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][52] ) );
  AOI22D2 U3258 ( .A1(n3412), .A2(\theRegs/managementDataOut[3][7] ), .B1(
        n3755), .B2(\theRegs/managementDataOut[2][7] ), .ZN(n2300) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[48].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[48].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][48] ) );
  AOI22D1 U3268 ( .A1(n3412), .A2(\theRegs/managementDataOut[3][5] ), .B1(
        n3755), .B2(\theRegs/managementDataOut[2][5] ), .ZN(n2292) );
  AOI22D2 U3273 ( .A1(n3412), .A2(\theRegs/managementDataOut[3][4] ), .B1(
        n3755), .B2(\theRegs/managementDataOut[2][4] ), .ZN(n2288) );
  NR2XD3 U4831 ( .A1(n3312), .A2(n3942), .ZN(n2243) );
  AOI22D2 U3278 ( .A1(n3412), .A2(\theRegs/managementDataOut[3][3] ), .B1(
        n3824), .B2(\theRegs/managementDataOut[2][3] ), .ZN(n2284) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][6] ) );
  CKND2 U3084 ( .I(n3887), .ZN(n3305) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][5] ) );
  AOI22D2 U3293 ( .A1(n3451), .A2(\theRegs/managementDataOut[3][0] ), .B1(
        n3824), .B2(\theRegs/managementDataOut[2][0] ), .ZN(n2272) );
  AOI22D2 U3288 ( .A1(n3451), .A2(\theRegs/managementDataOut[3][1] ), .B1(
        n3824), .B2(\theRegs/managementDataOut[2][1] ), .ZN(n2276) );
  AOI22D4 U3283 ( .A1(n3451), .A2(\theRegs/managementDataOut[3][2] ), .B1(
        n3824), .B2(\theRegs/managementDataOut[2][2] ), .ZN(n2280) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[64].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][64] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[2].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[2].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][2] ) );
  ND4D8 U2808 ( .A1(n3981), .A2(n3751), .A3(n3851), .A4(n3213), .ZN(n2183) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][6] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[9].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][9] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[28].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][28] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[9].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[9].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][9] ) );
  AOI22D4 U3263 ( .A1(n3451), .A2(\theRegs/managementDataOut[3][6] ), .B1(
        n3842), .B2(\theRegs/managementDataOut[2][6] ), .ZN(n2296) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[6].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[6].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][6] ) );
  AOI22D4 U3307 ( .A1(n3462), .A2(\theRegs/completionDataOut[6][67] ), .B1(
        n3909), .B2(\theRegs/completionDataOut[7][67] ), .ZN(n2575) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[27].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][27] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[24].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][24] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[27].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[27].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][27] ) );
  AOI22D4 U3308 ( .A1(n3569), .A2(\theRegs/completionDataOut[3][67] ), .B1(
        n3842), .B2(\theRegs/completionDataOut[2][67] ), .ZN(n2576) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[44].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[44].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][44] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[36].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][36] ) );
  AOI22D4 U3318 ( .A1(n3569), .A2(\theRegs/completionDataOut[3][65] ), .B1(
        n3842), .B2(\theRegs/completionDataOut[2][65] ), .ZN(n2568) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[29].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[29].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][29] ) );
  AO21D4 U2277 ( .A1(n3140), .A2(n3292), .B(n4117), .Z(n2232) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][4] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][8] ) );
  AOI22D4 U3313 ( .A1(n3569), .A2(\theRegs/completionDataOut[3][66] ), .B1(
        n3842), .B2(\theRegs/completionDataOut[2][66] ), .ZN(n2572) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][8] ) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[55].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][55] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[35].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][35] ) );
  BUFFD2 U3028 ( .I(n4038), .Z(n3294) );
  AOI22D4 U3317 ( .A1(n3462), .A2(\theRegs/completionDataOut[6][65] ), .B1(
        n3909), .B2(\theRegs/completionDataOut[7][65] ), .ZN(n2567) );
  AOI22D4 U3303 ( .A1(n3569), .A2(\theRegs/completionDataOut[3][68] ), .B1(
        n3916), .B2(\theRegs/completionDataOut[2][68] ), .ZN(n2580) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[55].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[55].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][55] ) );
  AOI22D4 U3320 ( .A1(n3505), .A2(\theRegs/completionDataOut[5][65] ), .B1(
        n3882), .B2(\theRegs/completionDataOut[4][65] ), .ZN(n2570) );
  BUFFD2 U4170 ( .I(n2202), .Z(n3311) );
  CKBD3 U4226 ( .I(n3940), .Z(n3336) );
  AOI22D4 U3253 ( .A1(\theRegs/managementDataOut[3][8] ), .A2(n3643), .B1(
        \theRegs/managementDataOut[2][8] ), .B2(n3916), .ZN(n2304) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[39].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[39].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][39] ) );
  AOI22D4 U3312 ( .A1(n3528), .A2(\theRegs/completionDataOut[6][66] ), .B1(
        n3909), .B2(\theRegs/completionDataOut[7][66] ), .ZN(n2571) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][0] ) );
  AOI22D4 U3315 ( .A1(n3932), .A2(\theRegs/completionDataOut[5][66] ), .B1(
        n3882), .B2(\theRegs/completionDataOut[4][66] ), .ZN(n2574) );
  AOI22D4 U3309 ( .A1(n3429), .A2(\theRegs/completionDataOut[1][67] ), .B1(
        n3801), .B2(\theRegs/completionDataOut[0][67] ), .ZN(n2577) );
  AOI22D4 U3270 ( .A1(n3932), .A2(\theRegs/managementDataOut[5][5] ), .B1(
        n3882), .B2(\theRegs/managementDataOut[4][5] ), .ZN(n2294) );
  AOI22D4 U3314 ( .A1(n3429), .A2(\theRegs/completionDataOut[1][66] ), .B1(
        n3931), .B2(\theRegs/completionDataOut[0][66] ), .ZN(n2573) );
  CKBD3 U2585 ( .I(decodeReadAddr2_i[0]), .Z(n3225) );
  AOI22D2 U3319 ( .A1(n3479), .A2(\theRegs/completionDataOut[1][65] ), .B1(
        n3931), .B2(\theRegs/completionDataOut[0][65] ), .ZN(n2569) );
  AOI22D4 U3299 ( .A1(n3479), .A2(\theRegs/completionDataOut[1][69] ), .B1(
        n3931), .B2(\theRegs/completionDataOut[0][69] ), .ZN(n2592) );
  AOI22D2 U3925 ( .A1(\theRegs/completionDataOut[2][7] ), .A2(n3881), .B1(
        \theRegs/completionDataOut[0][7] ), .B2(n3835), .ZN(n2830) );
  AO21D2 U2267 ( .A1(n3140), .A2(n3300), .B(reset_i), .Z(n2216) );
  AOI22D4 U3310 ( .A1(n3932), .A2(\theRegs/completionDataOut[5][67] ), .B1(
        n3882), .B2(\theRegs/completionDataOut[4][67] ), .ZN(n2578) );
  AOI22D2 U3910 ( .A1(\theRegs/completionDataOut[2][10] ), .A2(n3881), .B1(
        \theRegs/completionDataOut[0][10] ), .B2(n3835), .ZN(n2818) );
  ND2D3 U4829 ( .A1(n3284), .A2(n3887), .ZN(n2248) );
  AOI22D2 U4120 ( .A1(\theRegs/completionDataOut[2][3] ), .A2(n3881), .B1(
        \theRegs/completionDataOut[0][3] ), .B2(n3835), .ZN(n2846) );
  AOI22D2 U3675 ( .A1(\theRegs/completionDataOut[2][44] ), .A2(n3881), .B1(
        \theRegs/completionDataOut[0][44] ), .B2(n3835), .ZN(n2682) );
  DFQD2 \theRegs/eachManagementReg[1].managementReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[1][4] ) );
  ND4D8 U2600 ( .A1(n3212), .A2(n3981), .A3(n3751), .A4(n3851), .ZN(n2180) );
  DFQD2 \theRegs/eachManagementReg[1].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[1][5] ) );
  ND2D2 U4825 ( .A1(n3887), .A2(nextTail_o[0]), .ZN(n2247) );
  NR2D2 U4165 ( .A1(n2236), .A2(n3980), .ZN(n2196) );
  AO21D2 U2283 ( .A1(n3874), .A2(n3286), .B(n4117), .Z(n2229) );
  DFQD2 \theRegs/eachManagementReg[1].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[1][7] ) );
  DFQD2 \theRegs/eachManagementReg[4].managementReg/eachEnDff[7].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[7].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[4][7] ) );
  CKBD3 U4225 ( .I(n2197), .Z(n3335) );
  AOI22D2 U3634 ( .A1(n3813), .A2(\theRegs/completionDataOut[2][3] ), .B1(
        n3967), .B2(\theRegs/completionDataOut[1][3] ), .ZN(n2321) );
  AOI22D2 U3614 ( .A1(n3813), .A2(\theRegs/completionDataOut[2][7] ), .B1(
        n3967), .B2(\theRegs/completionDataOut[1][7] ), .ZN(n2337) );
  DFQD2 \theRegs/eachManagementReg[1].managementReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[1].managementReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[1][1] ) );
  NR3D4 U4205 ( .A1(n3229), .A2(n3226), .A3(n3228), .ZN(n3129) );
  DFQD2 \theRegs/eachManagementReg[5].managementReg/eachEnDff[3].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[5].managementReg/eachEnDff[3].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[5][3] ) );
  ND4D8 U3456 ( .A1(n2462), .A2(n2461), .A3(n2460), .A4(n2459), .ZN(
        commitReadData_o[38]) );
  ND4D8 U3626 ( .A1(n2326), .A2(n2325), .A3(n2324), .A4(n2323), .ZN(
        commitReadData_o[4]) );
  ND4D8 U3641 ( .A1(n2314), .A2(n2313), .A3(n2312), .A4(n2311), .ZN(
        commitReadData_o[1]) );
  CKBD4 U2914 ( .I(n2585), .Z(n3276) );
  BUFFD2 U3053 ( .I(n2584), .Z(n3300) );
  CKBD4 U3041 ( .I(n2583), .Z(n3298) );
  CKBD4 U2786 ( .I(n3129), .Z(n3251) );
  CKBD4 U2807 ( .I(n3128), .Z(n3259) );
  CKBD4 U2862 ( .I(n2860), .Z(n3265) );
  CKBD3 U3016 ( .I(n2587), .Z(n3292) );
  CKBD3 U3083 ( .I(\add_x_7/n1 ), .Z(n3304) );
  CKBD4 U2798 ( .I(n3129), .Z(n3252) );
  CKBD4 U2821 ( .I(n4006), .Z(n3260) );
  OAI32D4 U4846 ( .A1(n3241), .A2(n3250), .A3(n2256), .B1(n2253), .B2(n4011), 
        .ZN(n1405) );
  AO21D4 U2272 ( .A1(n3874), .A2(n3297), .B(n4117), .Z(n2212) );
  CKBD4 U3017 ( .I(n4038), .Z(n3293) );
  CKBD4 U2999 ( .I(n4008), .Z(n3289) );
  AOI22D4 U3282 ( .A1(n3374), .A2(\theRegs/managementDataOut[6][2] ), .B1(
        n3703), .B2(\theRegs/managementDataOut[7][2] ), .ZN(n2279) );
  AOI22D4 U3272 ( .A1(n3403), .A2(\theRegs/managementDataOut[6][4] ), .B1(
        n3829), .B2(\theRegs/managementDataOut[7][4] ), .ZN(n2287) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[31].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[31].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][31] ) );
  AOI22D4 U3267 ( .A1(n3452), .A2(\theRegs/managementDataOut[6][5] ), .B1(
        n3829), .B2(\theRegs/managementDataOut[7][5] ), .ZN(n2291) );
  CKBD3 U3100 ( .I(n2201), .Z(n3309) );
  AOI22D4 U3257 ( .A1(n3452), .A2(\theRegs/managementDataOut[6][7] ), .B1(
        n3829), .B2(\theRegs/managementDataOut[7][7] ), .ZN(n2299) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][1] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][4] ) );
  INR2XD1 U4828 ( .A1(n2243), .B1(n2248), .ZN(n2228) );
  AOI22D4 U3287 ( .A1(n3452), .A2(\theRegs/managementDataOut[6][1] ), .B1(
        n3829), .B2(\theRegs/managementDataOut[7][1] ), .ZN(n2275) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[61].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[61].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][61] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[64].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[64].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][64] ) );
  AOI22D4 U3277 ( .A1(n3452), .A2(\theRegs/managementDataOut[6][3] ), .B1(
        n3829), .B2(\theRegs/managementDataOut[7][3] ), .ZN(n2283) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[35].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[35].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][35] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[37].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[37].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][37] ) );
  NR2D2 U4179 ( .A1(n2247), .A2(n2220), .ZN(n2213) );
  DFQD2 \theRegs/eachCompletionReg[6].completionReg/eachEnDff[4].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[6].completionReg/eachEnDff[4].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[6][4] ) );
  AOI22D2 U3292 ( .A1(n3452), .A2(\theRegs/managementDataOut[6][0] ), .B1(
        n3968), .B2(\theRegs/managementDataOut[7][0] ), .ZN(n2271) );
  NR3D3 U4203 ( .A1(n3230), .A2(n3226), .A3(n3228), .ZN(n3133) );
  AOI22D2 U3467 ( .A1(n3461), .A2(\theRegs/completionDataOut[6][36] ), .B1(
        n3968), .B2(\theRegs/completionDataOut[7][36] ), .ZN(n2451) );
  AOI22D2 U3462 ( .A1(n3461), .A2(\theRegs/completionDataOut[6][37] ), .B1(
        n3968), .B2(\theRegs/completionDataOut[7][37] ), .ZN(n2455) );
  AOI22D2 U3622 ( .A1(n3461), .A2(\theRegs/completionDataOut[6][5] ), .B1(
        n3968), .B2(\theRegs/completionDataOut[7][5] ), .ZN(n2327) );
  NR3D3 U4202 ( .A1(n3225), .A2(n3230), .A3(n3228), .ZN(n3132) );
  AOI22D2 U3944 ( .A1(\theRegs/completionDataOut[3][30] ), .A2(n3837), .B1(
        \theRegs/completionDataOut[1][30] ), .B2(n3788), .ZN(n3010) );
  AOI22D2 U3959 ( .A1(\theRegs/completionDataOut[3][33] ), .A2(n3837), .B1(
        \theRegs/completionDataOut[1][33] ), .B2(n3788), .ZN(n2998) );
  INR2XD2 U2415 ( .A1(n2200), .B1(n2241), .ZN(n2202) );
  AOI22D2 U4014 ( .A1(\theRegs/completionDataOut[3][43] ), .A2(n3816), .B1(
        \theRegs/completionDataOut[1][43] ), .B2(n3769), .ZN(n2958) );
  AOI22D2 U3612 ( .A1(n3461), .A2(\theRegs/completionDataOut[6][7] ), .B1(
        n3968), .B2(\theRegs/completionDataOut[7][7] ), .ZN(n2335) );
  DFQD2 \theRegs/eachManagementReg[4].managementReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[4][5] ) );
  AOI22D4 U3106 ( .A1(n3513), .A2(\theRegs/completionDataOut[6][0] ), .B1(
        n3968), .B2(\theRegs/completionDataOut[7][0] ), .ZN(n2307) );
  CKND2 U2982 ( .I(n2207), .ZN(n3285) );
  DFQD2 \theRegs/eachManagementReg[2].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[2].managementReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[2][8] ) );
  DFQD2 \theRegs/eachManagementReg[4].managementReg/eachEnDff[8].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[4].managementReg/eachEnDff[8].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[4][8] ) );
  AOI21D4 U4819 ( .A1(n2268), .A2(\add_x_6/n1 ), .B(n3885), .ZN(n2210) );
  BUFFD2 U2260 ( .I(updateHead_i), .Z(n3140) );
  CKBD4 U2913 ( .I(n2585), .Z(n3275) );
  CKBD3 U2917 ( .I(n2856), .Z(n3279) );
  CKBD3 U2844 ( .I(n2855), .Z(n3263) );
  CKBD4 U2804 ( .I(n2859), .Z(n3257) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[49].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[49].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][49] ) );
  CKND2 U2597 ( .I(n3229), .ZN(n3230) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[22].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[22].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][22] ) );
  INR2XD1 U2666 ( .A1(n3791), .B1(n2232), .ZN(n2194) );
  NR2D2 U4162 ( .A1(n2212), .A2(n2180), .ZN(n2182) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[26].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][26] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[5].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[5].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][5] ) );
  CKBD3 U4207 ( .I(n2178), .Z(n3317) );
  CKBD3 U4191 ( .I(n2181), .Z(n3313) );
  AOI22D4 U3302 ( .A1(n3528), .A2(\theRegs/completionDataOut[6][68] ), .B1(
        n4010), .B2(\theRegs/completionDataOut[7][68] ), .ZN(n2579) );
  CKBD3 U4222 ( .I(n2179), .Z(n3332) );
  NR2D3 U4156 ( .A1(n2200), .A2(n2241), .ZN(n2201) );
  AOI22D2 U3627 ( .A1(n3513), .A2(\theRegs/completionDataOut[6][4] ), .B1(
        n4010), .B2(\theRegs/completionDataOut[7][4] ), .ZN(n2323) );
  NR2D2 U4161 ( .A1(n3976), .A2(n2223), .ZN(n2187) );
  AOI22D2 U3642 ( .A1(n3513), .A2(\theRegs/completionDataOut[6][1] ), .B1(
        n4010), .B2(\theRegs/completionDataOut[7][1] ), .ZN(n2311) );
  AOI22D2 U3109 ( .A1(n3882), .A2(\theRegs/completionDataOut[4][0] ), .B1(
        n3933), .B2(\theRegs/completionDataOut[0][0] ), .ZN(n2310) );
  AOI22D2 U3459 ( .A1(n3916), .A2(\theRegs/completionDataOut[2][38] ), .B1(
        n3479), .B2(\theRegs/completionDataOut[1][38] ), .ZN(n2461) );
  AOI22D2 U3473 ( .A1(n3932), .A2(\theRegs/completionDataOut[5][35] ), .B1(
        n3643), .B2(\theRegs/completionDataOut[3][35] ), .ZN(n2448) );
  AN3XD1 U2298 ( .A1(n3233), .A2(n3234), .A3(n3232), .Z(n2860) );
  CKBD4 U2901 ( .I(n2862), .Z(n3273) );
  CKBD3 U2915 ( .I(n3131), .Z(n3277) );
  CKBD3 U2824 ( .I(n3130), .Z(n3261) );
  CKBD4 U2936 ( .I(n2856), .Z(n3280) );
  CKBD4 U2866 ( .I(n3645), .Z(n3269) );
  CKBD4 U2845 ( .I(n3977), .Z(n3264) );
  BUFFD2 U2881 ( .I(n2858), .Z(n3271) );
  CKBD3 U2864 ( .I(n2861), .Z(n3267) );
  BUFFD2 U2652 ( .I(n3984), .Z(n3236) );
  BUFFD6 U2865 ( .I(n2861), .Z(n3268) );
  BUFFD6 U2902 ( .I(n2862), .Z(n3274) );
  CKBD4 U2916 ( .I(n3131), .Z(n3278) );
  CKBD4 U2841 ( .I(n3840), .Z(n3262) );
  CKBD4 U2898 ( .I(n2858), .Z(n3272) );
  CKBD4 U2655 ( .I(n3984), .Z(n3237) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[34].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[34].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][34] ) );
  OR2XD1 U2303 ( .A1(n3233), .A2(n3231), .Z(n2596) );
  INR2XD1 U2918 ( .A1(n3790), .B1(n2229), .ZN(n2191) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[24].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[24].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][24] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[26].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][26] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[47].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[47].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][47] ) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[57].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[57].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][57] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[36].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[36].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][36] ) );
  DFQD2 \theRegs/eachCompletionReg[3].completionReg/eachEnDff[1].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[3].completionReg/eachEnDff[1].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[3][1] ) );
  ND2D2 U4843 ( .A1(n3794), .A2(n2251), .ZN(n2256) );
  CKND4 U2595 ( .I(n3227), .ZN(n3228) );
  BUFFD2 U2632 ( .I(decodeReadAddr1_i[2]), .Z(n3234) );
  CKND2 U4187 ( .I(n2268), .ZN(n3312) );
  AOI221D4 U3005 ( .A1(n3793), .A2(n3983), .B1(n3312), .B2(n2262), .C(n2264), 
        .ZN(n1401) );
  BUFFD6 U2956 ( .I(n3135), .Z(n3282) );
  BUFFD6 U2878 ( .I(n3645), .Z(n3270) );
  AOI221D4 U3004 ( .A1(n3793), .A2(n3285), .B1(n3312), .B2(n2265), .C(n2264), 
        .ZN(n1400) );
  NR2D2 U4172 ( .A1(n2220), .A2(n4028), .ZN(n2217) );
  NR2D2 U4204 ( .A1(n3230), .A2(n2870), .ZN(n3131) );
  DFQD2 \theRegs/eachCompletionReg[0].completionReg/eachEnDff[30].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[0].completionReg/eachEnDff[30].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[0][30] ) );
  CKND2 U2633 ( .I(n3234), .ZN(n3235) );
  CKBD4 U2998 ( .I(n3688), .Z(n3288) );
  NR2XD1 U2293 ( .A1(n3234), .A2(n2596), .ZN(n2862) );
  CKND3 U2661 ( .I(tailReset), .ZN(n3239) );
  AOI22D2 U3643 ( .A1(n3718), .A2(\theRegs/completionDataOut[5][1] ), .B1(
        n3643), .B2(\theRegs/completionDataOut[3][1] ), .ZN(n2312) );
  NR2D2 U4163 ( .A1(n2232), .A2(n3978), .ZN(n2193) );
  NR2XD3 U4821 ( .A1(n3306), .A2(n2248), .ZN(\add_x_6/n1 ) );
  DFQD2 \theRegs/eachManagementReg[7].managementReg/eachEnDff[0].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachManagementReg[7].managementReg/eachEnDff[0].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/managementDataOut[7][0] ) );
  NR2D2 U4167 ( .A1(n2177), .A2(n2209), .ZN(n2178) );
  AOI22D2 U3674 ( .A1(\theRegs/completionDataOut[3][44] ), .A2(n3768), .B1(
        \theRegs/completionDataOut[1][44] ), .B2(n3815), .ZN(n2681) );
  NR2D3 U4171 ( .A1(n2217), .A2(n2216), .ZN(n2218) );
  DFQD2 \theRegs/eachCompletionReg[4].completionReg/eachEnDff[28].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[4].completionReg/eachEnDff[28].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[4][28] ) );
  NR2D3 U4126 ( .A1(n3235), .A2(n2596), .ZN(n2858) );
  NR2D2 U4199 ( .A1(n2598), .A2(n3235), .ZN(n2861) );
  ND2D1 U4198 ( .A1(n3226), .A2(n3228), .ZN(n2870) );
  NR2D3 U4189 ( .A1(n2229), .A2(n2228), .ZN(n2230) );
  NR2D2 U4166 ( .A1(n2229), .A2(n3979), .ZN(n2190) );
  AOI21D2 U4609 ( .A1(n3239), .A2(n3974), .B(n4031), .ZN(n1403) );
  CKBD4 U2997 ( .I(n3688), .Z(n3287) );
  NR2XD1 U4159 ( .A1(n4031), .A2(n2252), .ZN(n2251) );
  ND2D3 U4822 ( .A1(n2268), .A2(n3689), .ZN(n2220) );
  BUFFD2 U3052 ( .I(n2583), .Z(n3299) );
  CKBD3 U4208 ( .I(n2190), .Z(n3318) );
  NR2XD1 U4160 ( .A1(\headTailManager/headReset ), .A2(n2269), .ZN(n2252) );
  CKBD3 U2983 ( .I(n2588), .Z(n3286) );
  NR2D3 U4201 ( .A1(n2598), .A2(n2594), .ZN(n2856) );
  CKBD4 U4214 ( .I(n2193), .Z(n3324) );
  CKBD3 U4211 ( .I(n2196), .Z(n3321) );
  CKBD3 U4232 ( .I(n2188), .Z(n3342) );
  CKBD3 U3040 ( .I(n2589), .Z(n3297) );
  ND2D1 U2309 ( .A1(n3231), .A2(n3235), .ZN(n2594) );
  INR2XD1 U2499 ( .A1(n4029), .B1(n2223), .ZN(n2188) );
  ND2D2 U2311 ( .A1(n3233), .A2(n3231), .ZN(n2598) );
  CKBD4 U3039 ( .I(n2589), .Z(n3296) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[26].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[26].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][26] ) );
  DFQD2 \theRegs/eachCompletionReg[7].completionReg/eachEnDff[25].enDff/theFlop/q_reg  ( 
        .D(
        \theRegs/eachCompletionReg[7].completionReg/eachEnDff[25].enDff/theFlop/N3 ), .CP(clk_i), .Q(\theRegs/completionDataOut[7][25] ) );
  CKBD4 U3029 ( .I(n2589), .Z(n3295) );
  BUFFD2 U4210 ( .I(n2196), .Z(n3320) );
  AOI22D2 U3520 ( .A1(n3399), .A2(\theRegs/completionDataOut[4][26] ), .B1(
        n3547), .B2(\theRegs/completionDataOut[0][26] ), .ZN(n2414) );
  CKBD4 U3000 ( .I(n3495), .Z(n3290) );
  AOI22D4 U3517 ( .A1(n3516), .A2(\theRegs/completionDataOut[6][26] ), .B1(
        n3843), .B2(\theRegs/completionDataOut[7][26] ), .ZN(n2411) );
  AOI22D4 U3512 ( .A1(n3516), .A2(\theRegs/completionDataOut[6][27] ), .B1(
        n3302), .B2(\theRegs/completionDataOut[7][27] ), .ZN(n2415) );
  CKBD4 U4215 ( .I(n2193), .Z(n3325) );
  CKBD4 U4209 ( .I(n2190), .Z(n3319) );
  CKBD4 U2942 ( .I(n3135), .Z(n3281) );
  NR2XD1 U2317 ( .A1(n3229), .A2(n2870), .ZN(n3135) );
  CKBD3 U2596 ( .I(decodeReadAddr2_i[2]), .Z(n3229) );
  AOI221XD4 U4847 ( .A1(n3250), .A2(n4041), .B1(n4011), .B2(n4041), .C(
        head_o[3]), .ZN(head_o[2]) );
  NR4D4 U4173 ( .A1(n3887), .A2(nextTail_o[0]), .A3(n2220), .A4(n2216), .ZN(
        n2219) );
  BUFFD1 U2738 ( .I(n3134), .Z(n3645) );
  CKBD3 U4233 ( .I(n3346), .Z(n3343) );
  CKBD3 U4234 ( .I(n3299), .Z(n3344) );
  CKBD3 U4235 ( .I(n3348), .Z(n3345) );
  CKBD3 U4236 ( .I(n3281), .Z(n3346) );
  CKBD4 U4237 ( .I(n3353), .Z(n3347) );
  BUFFD2 U4238 ( .I(n3344), .Z(n3348) );
  CKBD4 U4239 ( .I(n3324), .Z(n3349) );
  CKBD3 U4240 ( .I(n3386), .Z(n3350) );
  CKBD3 U4241 ( .I(n3361), .Z(n3351) );
  CKBD3 U4242 ( .I(n3300), .Z(n3352) );
  CKBD3 U4243 ( .I(n3346), .Z(n3353) );
  CKBD4 U4244 ( .I(n3348), .Z(n3354) );
  CKBD3 U4245 ( .I(n3371), .Z(n3355) );
  CKBD3 U4246 ( .I(n3385), .Z(n3356) );
  CKBD3 U4247 ( .I(n3321), .Z(n3357) );
  CKBD3 U4248 ( .I(n3368), .Z(n3358) );
  CKBD4 U4249 ( .I(n3369), .Z(n3359) );
  CKBD3 U4250 ( .I(n3318), .Z(n3360) );
  BUFFD2 U4251 ( .I(n3324), .Z(n3361) );
  CKBD4 U4252 ( .I(n3352), .Z(n3362) );
  CKBD3 U4253 ( .I(n3296), .Z(n3363) );
  CKBD3 U4254 ( .I(n3381), .Z(n3364) );
  CKBD3 U4257 ( .I(n3384), .Z(n3365) );
  CKBD3 U4258 ( .I(n3517), .Z(n3366) );
  CKBD3 U4259 ( .I(n3382), .Z(n3367) );
  CKBD4 U4260 ( .I(n3353), .Z(n3368) );
  CKBD3 U4261 ( .I(n3354), .Z(n3369) );
  CKBD3 U4262 ( .I(n3363), .Z(n3370) );
  BUFFD2 U4263 ( .I(n3290), .Z(n3371) );
  BUFFD0 U4264 ( .I(n2195), .Z(n3372) );
  BUFFD1 U4265 ( .I(n3399), .Z(n3373) );
  CKBD3 U4266 ( .I(n3403), .Z(n3374) );
  CKBD3 U4267 ( .I(n3404), .Z(n3375) );
  CKBD3 U4268 ( .I(n3425), .Z(n3376) );
  CKBD3 U4269 ( .I(n3400), .Z(n3377) );
  CKBD4 U4270 ( .I(n3286), .Z(n3378) );
  CKBD4 U4271 ( .I(n3261), .Z(n3379) );
  CKBD4 U4272 ( .I(n3323), .Z(n3380) );
  BUFFD2 U4273 ( .I(n3324), .Z(n3381) );
  CKBD3 U4274 ( .I(n3318), .Z(n3382) );
  CKBD4 U4275 ( .I(n3371), .Z(n3383) );
  BUFFD2 U4276 ( .I(n3321), .Z(n3384) );
  BUFFD2 U4277 ( .I(n3276), .Z(n3385) );
  BUFFD2 U4278 ( .I(n3287), .Z(n3386) );
  CKBD4 U4279 ( .I(n3342), .Z(n3387) );
  CKBD3 U4280 ( .I(n3417), .Z(n3388) );
  CKBD3 U4281 ( .I(n3420), .Z(n3389) );
  CKBD3 U4282 ( .I(n3421), .Z(n3390) );
  CKBD3 U4283 ( .I(n3423), .Z(n3391) );
  BUFFD1 U4284 ( .I(n3491), .Z(n3392) );
  BUFFD2 U4285 ( .I(n3320), .Z(n3393) );
  CKBD3 U4286 ( .I(n3236), .Z(n3394) );
  CKBD3 U4287 ( .I(n3418), .Z(n3395) );
  CKBD3 U4288 ( .I(n3419), .Z(n3396) );
  CKBD3 U4289 ( .I(n3267), .Z(n3397) );
  CKBD4 U4290 ( .I(n3277), .Z(n3398) );
  CKBD4 U4291 ( .I(n3369), .Z(n3399) );
  CKBD4 U4292 ( .I(n3370), .Z(n3400) );
  CKBD3 U4293 ( .I(n3342), .Z(n3401) );
  CKBD4 U4294 ( .I(n3378), .Z(n3402) );
  BUFFD2 U4295 ( .I(n3297), .Z(n3403) );
  BUFFD2 U4296 ( .I(n3368), .Z(n3404) );
  CKBD3 U4297 ( .I(n3449), .Z(n3405) );
  CKBD3 U4298 ( .I(n3488), .Z(n3406) );
  BUFFD1 U4299 ( .I(n3490), .Z(n3407) );
  CKBD3 U4300 ( .I(n3262), .Z(n3408) );
  CKBD3 U4301 ( .I(n3271), .Z(n3409) );
  CKBD3 U4302 ( .I(n3263), .Z(n3410) );
  CKBD3 U4303 ( .I(n3275), .Z(n3411) );
  BUFFD2 U4304 ( .I(n3451), .Z(n3412) );
  CKBD3 U4305 ( .I(n3453), .Z(n3413) );
  CKBD3 U4306 ( .I(n3265), .Z(n3414) );
  CKBD4 U4307 ( .I(n3270), .Z(n3415) );
  CKBD3 U4308 ( .I(n3273), .Z(n3416) );
  BUFFD2 U4309 ( .I(n3324), .Z(n3417) );
  CKBD3 U4310 ( .I(n3318), .Z(n3418) );
  CKBD4 U4311 ( .I(n3383), .Z(n3419) );
  BUFFD2 U4312 ( .I(n3357), .Z(n3420) );
  BUFFD1 U4313 ( .I(n3386), .Z(n3421) );
  CKBD4 U4314 ( .I(n3385), .Z(n3422) );
  CKBD3 U4315 ( .I(n3323), .Z(n3423) );
  CKBD4 U4316 ( .I(n3398), .Z(n3424) );
  BUFFD1 U4317 ( .I(n3332), .Z(n3425) );
  CKBD3 U4318 ( .I(n3450), .Z(n3426) );
  CKBD3 U4319 ( .I(n3477), .Z(n3427) );
  BUFFD1 U4320 ( .I(n3478), .Z(n3428) );
  CKBD3 U4321 ( .I(n3479), .Z(n3429) );
  BUFFD1 U4322 ( .I(n3480), .Z(n3430) );
  CKBD3 U4323 ( .I(n3481), .Z(n3431) );
  BUFFD2 U4324 ( .I(n3482), .Z(n3432) );
  BUFFD2 U4325 ( .I(n3483), .Z(n3433) );
  CKBD3 U4326 ( .I(n3486), .Z(n3434) );
  CKBD3 U4327 ( .I(n3549), .Z(n3435) );
  CKBD3 U4328 ( .I(n3555), .Z(n3436) );
  CKBD3 U4329 ( .I(n3561), .Z(n3437) );
  BUFFD1 U4330 ( .I(n3563), .Z(n3438) );
  BUFFD2 U4331 ( .I(n3278), .Z(n3439) );
  CKBD3 U4332 ( .I(n3257), .Z(n3440) );
  CKBD3 U4333 ( .I(n3279), .Z(n3441) );
  CKBD3 U4334 ( .I(n3489), .Z(n3442) );
  CKBD3 U4335 ( .I(n3255), .Z(n3443) );
  CKBD3 U4336 ( .I(n3518), .Z(n3444) );
  CKBD4 U4337 ( .I(n3264), .Z(n3445) );
  CKBD3 U4338 ( .I(n3521), .Z(n3446) );
  CKBD4 U4339 ( .I(n3282), .Z(n3447) );
  CKBD3 U4340 ( .I(n3309), .Z(n3448) );
  BUFFD2 U4341 ( .I(n3400), .Z(n3449) );
  CKBD3 U4342 ( .I(n3342), .Z(n3450) );
  CKBD3 U4343 ( .I(n3402), .Z(n3451) );
  CKBD4 U4344 ( .I(n3403), .Z(n3452) );
  BUFFD2 U4345 ( .I(n3320), .Z(n3453) );
  CKBD4 U4346 ( .I(n3379), .Z(n3454) );
  CKBD4 U4347 ( .I(n3416), .Z(n3455) );
  CKBD4 U4348 ( .I(n3411), .Z(n3456) );
  CKBD3 U4349 ( .I(n3295), .Z(n3457) );
  CKBD4 U4350 ( .I(n3272), .Z(n3458) );
  CKBD4 U4351 ( .I(n3274), .Z(n3459) );
  CKBD3 U4352 ( .I(n3512), .Z(n3460) );
  CKBD3 U4353 ( .I(n3513), .Z(n3461) );
  CKBD3 U4354 ( .I(n3528), .Z(n3462) );
  CKBD3 U4355 ( .I(n3550), .Z(n3463) );
  CKBD3 U4356 ( .I(n3523), .Z(n3464) );
  CKBD3 U4357 ( .I(n3554), .Z(n3465) );
  BUFFD2 U4358 ( .I(n3560), .Z(n3466) );
  CKBD3 U4359 ( .I(n3514), .Z(n3467) );
  CKBD3 U4360 ( .I(n3520), .Z(n3468) );
  CKBD3 U4361 ( .I(n3553), .Z(n3469) );
  CKBD3 U4362 ( .I(n3556), .Z(n3470) );
  CKBD4 U4363 ( .I(n3280), .Z(n3471) );
  CKBD3 U4364 ( .I(n3291), .Z(n3472) );
  BUFFD2 U4365 ( .I(n3326), .Z(n3473) );
  CKBD3 U4366 ( .I(n3558), .Z(n3474) );
  CKBD3 U4367 ( .I(n3311), .Z(n3475) );
  CKBD3 U4368 ( .I(n3253), .Z(n3476) );
  BUFFD2 U4369 ( .I(n3324), .Z(n3477) );
  CKBD3 U4370 ( .I(n3318), .Z(n3478) );
  BUFFD2 U4371 ( .I(n3419), .Z(n3479) );
  CKBD4 U4372 ( .I(n3321), .Z(n3480) );
  BUFFD2 U4373 ( .I(n3421), .Z(n3481) );
  CKBD3 U4374 ( .I(n3422), .Z(n3482) );
  CKBD3 U4375 ( .I(n3323), .Z(n3483) );
  CKBD3 U4376 ( .I(n3393), .Z(n3484) );
  CKBD4 U4377 ( .I(n3458), .Z(n3485) );
  BUFFD2 U4378 ( .I(n3414), .Z(n3486) );
  CKBD4 U4379 ( .I(n3397), .Z(n3487) );
  CKBD3 U4380 ( .I(n3394), .Z(n3488) );
  CKBD4 U4381 ( .I(n3259), .Z(n3489) );
  CKBD4 U4382 ( .I(n3268), .Z(n3490) );
  CKBD3 U4383 ( .I(n3317), .Z(n3491) );
  CKBD4 U4384 ( .I(n3410), .Z(n3492) );
  CKBD4 U4385 ( .I(n3515), .Z(n3493) );
  CKBD4 U4386 ( .I(n3516), .Z(n3494) );
  BUFFD1 U4387 ( .I(n2586), .Z(n3495) );
  CKBD3 U4388 ( .I(n3593), .Z(n3496) );
  CKBD3 U4389 ( .I(n3594), .Z(n3497) );
  CKBD3 U4390 ( .I(n3635), .Z(n3498) );
  BUFFD1 U4391 ( .I(n3638), .Z(n3499) );
  BUFFD2 U4392 ( .I(n3641), .Z(n3500) );
  CKBD3 U4393 ( .I(n3562), .Z(n3501) );
  CKBD3 U4394 ( .I(n3596), .Z(n3502) );
  CKBD3 U4395 ( .I(n3603), .Z(n3503) );
  CKBD3 U4396 ( .I(n3685), .Z(n3504) );
  CKBD3 U4397 ( .I(n3932), .Z(n3505) );
  CKBD3 U4398 ( .I(n3548), .Z(n3506) );
  CKBD4 U4399 ( .I(n3551), .Z(n3507) );
  CKBD4 U4400 ( .I(n3595), .Z(n3508) );
  CKBD3 U4401 ( .I(n3599), .Z(n3509) );
  CKBD3 U4402 ( .I(n3546), .Z(n3510) );
  CKBD3 U4403 ( .I(n3547), .Z(n3511) );
  CKBD3 U4404 ( .I(n3342), .Z(n3512) );
  CKBD3 U4405 ( .I(n3452), .Z(n3513) );
  CKBD3 U4406 ( .I(n3454), .Z(n3514) );
  CKBD4 U4407 ( .I(n3456), .Z(n3515) );
  CKBD4 U4408 ( .I(n3457), .Z(n3516) );
  CKBD4 U4409 ( .I(n3362), .Z(n3517) );
  CKBD4 U4410 ( .I(n3415), .Z(n3518) );
  CKBD4 U4411 ( .I(n3488), .Z(n3519) );
  CKBD3 U4412 ( .I(n3309), .Z(n3520) );
  CKBD3 U4413 ( .I(n3408), .Z(n3521) );
  CKBD4 U4414 ( .I(n3476), .Z(n3522) );
  CKBD3 U4415 ( .I(n3269), .Z(n3523) );
  CKBD4 U4416 ( .I(n3440), .Z(n3524) );
  CKBD4 U4417 ( .I(n3441), .Z(n3525) );
  CKBD4 U4418 ( .I(n3237), .Z(n3526) );
  CKBD4 U4419 ( .I(n3256), .Z(n3527) );
  BUFFD2 U4420 ( .I(n3449), .Z(n3528) );
  CKBD3 U4421 ( .I(n3590), .Z(n3529) );
  CKBD3 U4422 ( .I(n3591), .Z(n3530) );
  CKBD3 U4423 ( .I(n3626), .Z(n3531) );
  CKBD3 U4424 ( .I(n3629), .Z(n3532) );
  CKBD3 U4425 ( .I(n3636), .Z(n3533) );
  CKBD3 U4426 ( .I(n3668), .Z(n3534) );
  BUFFD1 U4427 ( .I(n3686), .Z(n3535) );
  CKBD3 U4428 ( .I(n3602), .Z(n3536) );
  CKBD3 U4429 ( .I(n3637), .Z(n3537) );
  CKBD3 U4430 ( .I(n3260), .Z(n3538) );
  BUFFD2 U4431 ( .I(n3589), .Z(n3539) );
  CKBD4 U4432 ( .I(n3592), .Z(n3540) );
  CKBD3 U4433 ( .I(n3628), .Z(n3541) );
  CKBD3 U4434 ( .I(n3630), .Z(n3542) );
  CKBD3 U4435 ( .I(n3631), .Z(n3543) );
  CKBD4 U4436 ( .I(n3633), .Z(n3544) );
  CKBD4 U4437 ( .I(n3288), .Z(n3545) );
  CKBD3 U4438 ( .I(n3321), .Z(n3546) );
  CKBD4 U4439 ( .I(n3482), .Z(n3547) );
  BUFFD2 U4440 ( .I(n3393), .Z(n3548) );
  BUFFD2 U4441 ( .I(n3424), .Z(n3549) );
  BUFFD2 U4442 ( .I(n3455), .Z(n3550) );
  CKBD3 U4443 ( .I(n3489), .Z(n3551) );
  CKBD4 U4444 ( .I(n3522), .Z(n3552) );
  CKBD4 U4445 ( .I(n3447), .Z(n3553) );
  CKBD4 U4446 ( .I(n3459), .Z(n3554) );
  CKBD3 U4447 ( .I(n3332), .Z(n3555) );
  CKBD4 U4448 ( .I(n3445), .Z(n3556) );
  CKBD4 U4449 ( .I(n3526), .Z(n3557) );
  CKBD3 U4450 ( .I(n3439), .Z(n3558) );
  CKBD3 U4451 ( .I(n3311), .Z(n3559) );
  CKBD4 U4452 ( .I(n3882), .Z(n3560) );
  CKBD3 U4453 ( .I(n3409), .Z(n3561) );
  BUFFD2 U4454 ( .I(n3293), .Z(n3562) );
  BUFFD2 U4455 ( .I(n3313), .Z(n3563) );
  CKBD4 U4456 ( .I(n3254), .Z(n3564) );
  CKBD4 U4457 ( .I(n3258), .Z(n3565) );
  CKBD3 U4458 ( .I(n3331), .Z(n3566) );
  BUFFD1 U4459 ( .I(n3627), .Z(n3567) );
  CKBD3 U4460 ( .I(n3634), .Z(n3568) );
  CKBD3 U4461 ( .I(n3643), .Z(n3569) );
  CKBD3 U4462 ( .I(n3673), .Z(n3570) );
  CKBD3 U4463 ( .I(n3676), .Z(n3571) );
  BUFFD2 U4464 ( .I(n3722), .Z(n3572) );
  CKBD3 U4465 ( .I(n3819), .Z(n3573) );
  CKBD3 U4466 ( .I(n3319), .Z(n3574) );
  CKBD3 U4467 ( .I(n3640), .Z(n3575) );
  CKBD3 U4468 ( .I(n3680), .Z(n3576) );
  CKBD3 U4469 ( .I(n3681), .Z(n3577) );
  CKBD3 U4470 ( .I(n3252), .Z(n3578) );
  CKBD3 U4471 ( .I(n3644), .Z(n3579) );
  CKBD3 U4472 ( .I(n3666), .Z(n3580) );
  CKBD3 U4473 ( .I(n3667), .Z(n3581) );
  CKBD3 U4474 ( .I(n3671), .Z(n3582) );
  CKBD3 U4475 ( .I(n3672), .Z(n3583) );
  CKBD3 U4476 ( .I(n3674), .Z(n3584) );
  CKBD3 U4477 ( .I(n3675), .Z(n3585) );
  CKBD3 U4478 ( .I(n3677), .Z(n3586) );
  CKBD3 U4479 ( .I(n3340), .Z(n3587) );
  BUFFD2 U4480 ( .I(n3308), .Z(n3588) );
  CKBD3 U4481 ( .I(n3342), .Z(n3589) );
  BUFFD2 U4482 ( .I(n3318), .Z(n3590) );
  BUFFD2 U4483 ( .I(n3481), .Z(n3591) );
  CKBD3 U4484 ( .I(n3523), .Z(n3592) );
  BUFFD2 U4485 ( .I(n3486), .Z(n3593) );
  BUFFD2 U4486 ( .I(n3487), .Z(n3594) );
  CKBD4 U4487 ( .I(n3492), .Z(n3595) );
  CKBD4 U4488 ( .I(n3490), .Z(n3596) );
  CKBD4 U4489 ( .I(n3560), .Z(n3597) );
  CKBD4 U4490 ( .I(n3561), .Z(n3598) );
  CKBD4 U4491 ( .I(n3471), .Z(n3599) );
  BUFFD2 U4492 ( .I(n3313), .Z(n3600) );
  CKBD4 U4493 ( .I(n3545), .Z(n3601) );
  CKBD4 U4494 ( .I(n3632), .Z(n3602) );
  CKBD4 U4495 ( .I(n3251), .Z(n3603) );
  CKBD4 U4496 ( .I(n3443), .Z(n3604) );
  CKBD4 U4497 ( .I(n3266), .Z(n3605) );
  BUFFD1 U4498 ( .I(n3665), .Z(n3606) );
  CKBD3 U4499 ( .I(n3683), .Z(n3607) );
  CKBD3 U4500 ( .I(n3719), .Z(n3608) );
  CKBD3 U4501 ( .I(n3733), .Z(n3609) );
  BUFFD1 U4502 ( .I(n3782), .Z(n3610) );
  CKBD3 U4503 ( .I(n3726), .Z(n3611) );
  CKBD3 U4504 ( .I(n3732), .Z(n3612) );
  CKBD3 U4505 ( .I(n3292), .Z(n3613) );
  CKBD3 U4506 ( .I(n3669), .Z(n3614) );
  CKBD3 U4507 ( .I(n3670), .Z(n3615) );
  CKBD3 U4508 ( .I(n3678), .Z(n3616) );
  CKBD3 U4509 ( .I(n3715), .Z(n3617) );
  CKBD3 U4510 ( .I(n3716), .Z(n3618) );
  CKBD3 U4511 ( .I(n3717), .Z(n3619) );
  CKBD3 U4512 ( .I(n3720), .Z(n3620) );
  CKBD4 U4513 ( .I(n3723), .Z(n3621) );
  CKBD3 U4514 ( .I(n3727), .Z(n3622) );
  CKBD3 U4515 ( .I(n3774), .Z(n3623) );
  CKBD3 U4516 ( .I(n3319), .Z(n3624) );
  CKBD4 U4517 ( .I(n3304), .Z(n3625) );
  BUFFD2 U4518 ( .I(n3514), .Z(n3626) );
  CKBD3 U4519 ( .I(n3323), .Z(n3627) );
  CKBD3 U4520 ( .I(n3309), .Z(n3628) );
  CKBD3 U4521 ( .I(n3518), .Z(n3629) );
  CKBD4 U4522 ( .I(n3485), .Z(n3630) );
  CKBD4 U4523 ( .I(n3521), .Z(n3631) );
  CKBD4 U4524 ( .I(n3331), .Z(n3632) );
  CKBD4 U4525 ( .I(n3525), .Z(n3633) );
  BUFFD2 U4526 ( .I(n3562), .Z(n3634) );
  CKBD3 U4527 ( .I(n3317), .Z(n3635) );
  BUFFD2 U4528 ( .I(n3524), .Z(n3636) );
  CKBD3 U4529 ( .I(n3527), .Z(n3637) );
  BUFFD2 U4530 ( .I(n3326), .Z(n3638) );
  CKBD4 U4531 ( .I(n3538), .Z(n3639) );
  BUFFD1 U4532 ( .I(n3322), .Z(n3640) );
  CKBD4 U4533 ( .I(n3301), .Z(n3641) );
  CKBD3 U4534 ( .I(n3302), .Z(n3642) );
  CKBD3 U4535 ( .I(n3451), .Z(n3643) );
  BUFFD2 U4536 ( .I(n3399), .Z(n3644) );
  BUFFD2 U4537 ( .I(n3718), .Z(n3646) );
  CKBD3 U4538 ( .I(n3721), .Z(n3647) );
  CKBD3 U4539 ( .I(n3766), .Z(n3648) );
  CKBD3 U4540 ( .I(n3767), .Z(n3649) );
  CKBD3 U4541 ( .I(n3768), .Z(n3650) );
  CKBD3 U4542 ( .I(n3769), .Z(n3651) );
  CKBD3 U4543 ( .I(n3775), .Z(n3652) );
  CKBD3 U4544 ( .I(n3776), .Z(n3653) );
  CKBD3 U4545 ( .I(n3778), .Z(n3654) );
  CKBD3 U4546 ( .I(n3788), .Z(n3655) );
  CKBD3 U4547 ( .I(n3725), .Z(n3656) );
  CKBD3 U4548 ( .I(n3787), .Z(n3657) );
  CKBD3 U4549 ( .I(n3714), .Z(n3658) );
  CKBD3 U4550 ( .I(n3773), .Z(n3659) );
  CKBD4 U4551 ( .I(n3779), .Z(n3660) );
  CKBD3 U4552 ( .I(n3724), .Z(n3661) );
  CKBD3 U4553 ( .I(n3730), .Z(n3662) );
  CKBD3 U4554 ( .I(n3781), .Z(n3663) );
  CKBD3 U4555 ( .I(n3289), .Z(n3664) );
  CKBD4 U4556 ( .I(n3321), .Z(n3665) );
  CKBD4 U4557 ( .I(n3549), .Z(n3666) );
  CKBD4 U4558 ( .I(n3550), .Z(n3667) );
  CKBD4 U4559 ( .I(n3515), .Z(n3668) );
  CKBD4 U4560 ( .I(n3551), .Z(n3669) );
  CKBD4 U4561 ( .I(n3595), .Z(n3670) );
  CKBD3 U4562 ( .I(n3519), .Z(n3671) );
  CKBD4 U4563 ( .I(n3556), .Z(n3672) );
  CKBD3 U4564 ( .I(n3553), .Z(n3673) );
  CKBD4 U4565 ( .I(n3557), .Z(n3674) );
  CKBD4 U4566 ( .I(n3558), .Z(n3675) );
  CKBD4 U4567 ( .I(n3554), .Z(n3676) );
  BUFFD2 U4568 ( .I(n3311), .Z(n3677) );
  CKBD4 U4569 ( .I(n3604), .Z(n3678) );
  CKBD3 U4570 ( .I(n3473), .Z(n3679) );
  CKBD3 U4571 ( .I(n3564), .Z(n3680) );
  CKBD3 U4572 ( .I(n3565), .Z(n3681) );
  CKBD4 U4573 ( .I(n3641), .Z(n3682) );
  BUFFD2 U4574 ( .I(n3472), .Z(n3683) );
  CKBD4 U4575 ( .I(n3578), .Z(n3684) );
  BUFFD2 U4576 ( .I(n3316), .Z(n3685) );
  CKBD4 U4577 ( .I(n3324), .Z(n3686) );
  CKBD4 U4578 ( .I(n3338), .Z(n3687) );
  BUFFD1 U4579 ( .I(n2588), .Z(n3688) );
  BUFFD1 U4580 ( .I(n2227), .Z(n3689) );
  BUFFD1 U4581 ( .I(n2210), .Z(n3690) );
  CKBD3 U4582 ( .I(n3814), .Z(n3691) );
  CKBD3 U4583 ( .I(n3815), .Z(n3692) );
  CKBD3 U4584 ( .I(n3816), .Z(n3693) );
  CKBD3 U4585 ( .I(n3817), .Z(n3694) );
  CKBD3 U4586 ( .I(n3821), .Z(n3695) );
  CKBD3 U4587 ( .I(n3822), .Z(n3696) );
  BUFFD2 U4588 ( .I(n3835), .Z(n3697) );
  CKBD3 U4589 ( .I(n3837), .Z(n3698) );
  CKBD3 U4590 ( .I(n3838), .Z(n3699) );
  BUFFD2 U4591 ( .I(n3784), .Z(n3700) );
  CKBD3 U4592 ( .I(n3785), .Z(n3701) );
  CKBD3 U4593 ( .I(n3786), .Z(n3702) );
  CKBD3 U4594 ( .I(head_o[3]), .Z(n3703) );
  CKBD3 U4595 ( .I(n3770), .Z(n3704) );
  CKBD3 U4596 ( .I(n3772), .Z(n3705) );
  CKBD3 U4597 ( .I(n3783), .Z(n3706) );
  CKBD4 U4598 ( .I(n3820), .Z(n3707) );
  CKBD4 U4599 ( .I(n3823), .Z(n3708) );
  CKBD3 U4600 ( .I(n3915), .Z(n3709) );
  CKBD3 U4601 ( .I(n3328), .Z(n3710) );
  CKBD3 U4602 ( .I(n3812), .Z(n3711) );
  CKBD4 U4603 ( .I(n3834), .Z(n3712) );
  CKBD3 U4604 ( .I(n3330), .Z(n3713) );
  CKBD4 U4605 ( .I(n3592), .Z(n3714) );
  CKBD4 U4606 ( .I(n3593), .Z(n3715) );
  CKBD4 U4607 ( .I(n3594), .Z(n3716) );
  CKBD3 U4608 ( .I(n3598), .Z(n3717) );
  CKBD4 U4610 ( .I(n3517), .Z(n3718) );
  CKBD4 U4611 ( .I(n3596), .Z(n3719) );
  CKBD4 U4612 ( .I(n3599), .Z(n3720) );
  BUFFD2 U4613 ( .I(n3634), .Z(n3721) );
  CKBD3 U4614 ( .I(n3332), .Z(n3722) );
  CKBD3 U4615 ( .I(n3603), .Z(n3723) );
  CKBD4 U4616 ( .I(n3625), .Z(n3724) );
  BUFFD2 U4617 ( .I(n3642), .Z(n3725) );
  CKBD3 U4618 ( .I(n3605), .Z(n3726) );
  BUFFD2 U4619 ( .I(n3308), .Z(n3727) );
  BUFFD2 U4620 ( .I(n3325), .Z(n3728) );
  CKBD4 U4621 ( .I(n3338), .Z(n3729) );
  CKBD3 U4622 ( .I(n3334), .Z(n3730) );
  CKBD4 U4623 ( .I(n3613), .Z(n3731) );
  BUFFD2 U4624 ( .I(n3341), .Z(n3732) );
  CKBD3 U4625 ( .I(n3298), .Z(n3733) );
  CKBD4 U4626 ( .I(n3771), .Z(n3734) );
  CKBD4 U4627 ( .I(n3777), .Z(n3735) );
  BUFFD1 U4628 ( .I(n3736), .Z(n2855) );
  CKBD3 U4629 ( .I(n3813), .Z(n3737) );
  BUFFD1 U4630 ( .I(n3836), .Z(n3738) );
  CKBD3 U4631 ( .I(n3861), .Z(n3739) );
  CKBD3 U4632 ( .I(n3862), .Z(n3740) );
  CKBD3 U4633 ( .I(n3866), .Z(n3741) );
  CKBD3 U4634 ( .I(n3868), .Z(n3742) );
  BUFFD1 U4635 ( .I(n3873), .Z(n3743) );
  CKBD3 U4637 ( .I(n3877), .Z(n3744) );
  BUFFD1 U4638 ( .I(n3879), .Z(n3745) );
  BUFFD2 U4639 ( .I(n3881), .Z(n3746) );
  CKBD3 U4640 ( .I(n3928), .Z(n3747) );
  BUFFD1 U4641 ( .I(n3333), .Z(n3748) );
  CKBD3 U4642 ( .I(n3827), .Z(n3749) );
  CKBD3 U4643 ( .I(n3933), .Z(n3750) );
  BUFFD2 U4644 ( .I(n3214), .Z(n3751) );
  BUFFD1 U4645 ( .I(n2230), .Z(n3752) );
  BUFFD1 U4646 ( .I(n2218), .Z(n3753) );
  CKBD3 U4647 ( .I(n3818), .Z(n3754) );
  BUFFD2 U4648 ( .I(n3824), .Z(n3755) );
  CKBD3 U4649 ( .I(n3863), .Z(n3756) );
  CKBD3 U4650 ( .I(n3864), .Z(n3757) );
  CKBD3 U4651 ( .I(n3867), .Z(n3758) );
  CKBD3 U4652 ( .I(n3870), .Z(n3759) );
  BUFFD2 U4653 ( .I(n3871), .Z(n3760) );
  CKBD3 U4654 ( .I(n3919), .Z(n3761) );
  BUFFD1 U4655 ( .I(n2210), .Z(n3762) );
  CKBD3 U4656 ( .I(n3828), .Z(n3763) );
  CKBD4 U4657 ( .I(n3860), .Z(n3764) );
  CKBD4 U4658 ( .I(n3878), .Z(n3765) );
  CKBD3 U4659 ( .I(n3309), .Z(n3766) );
  CKBD4 U4660 ( .I(n3629), .Z(n3767) );
  CKBD3 U4661 ( .I(n3630), .Z(n3768) );
  CKBD3 U4662 ( .I(n3631), .Z(n3769) );
  CKBD4 U4663 ( .I(n3678), .Z(n3770) );
  CKBD4 U4664 ( .I(n3597), .Z(n3771) );
  CKBD4 U4665 ( .I(n3633), .Z(n3772) );
  CKBD4 U4666 ( .I(n3636), .Z(n3773) );
  BUFFD2 U4667 ( .I(n3313), .Z(n3774) );
  CKBD3 U4668 ( .I(n3317), .Z(n3775) );
  CKBD3 U4669 ( .I(n3637), .Z(n3776) );
  CKBD4 U4670 ( .I(n3316), .Z(n3777) );
  CKBD3 U4671 ( .I(n3601), .Z(n3778) );
  CKBD3 U4672 ( .I(n3639), .Z(n3779) );
  CKBD3 U4673 ( .I(n3330), .Z(n3780) );
  BUFFD2 U4674 ( .I(n3310), .Z(n3781) );
  BUFFD2 U4675 ( .I(n3340), .Z(n3782) );
  CKBD3 U4676 ( .I(n3336), .Z(n3783) );
  CKBD3 U4677 ( .I(n3811), .Z(n3784) );
  CKBD3 U4678 ( .I(n3339), .Z(n3785) );
  BUFFD1 U4679 ( .I(n3337), .Z(n3786) );
  BUFFD2 U4680 ( .I(n3329), .Z(n3787) );
  CKBD3 U4681 ( .I(n3626), .Z(n3788) );
  BUFFD0 U4682 ( .I(n2855), .Z(n3789) );
  BUFFD0 U4683 ( .I(n2189), .Z(n3790) );
  BUFFD0 U4684 ( .I(n2192), .Z(n3791) );
  BUFFD1 U4685 ( .I(n2227), .Z(n3792) );
  BUFFD1 U4686 ( .I(n2268), .Z(n3793) );
  BUFFD1 U4687 ( .I(n3874), .Z(n3794) );
  CKBD3 U4688 ( .I(n3880), .Z(n3795) );
  CKBD3 U4689 ( .I(n3907), .Z(n3796) );
  CKBD3 U4690 ( .I(n3911), .Z(n3797) );
  CKBD3 U4691 ( .I(n3913), .Z(n3798) );
  CKBD3 U4692 ( .I(n3929), .Z(n3799) );
  BUFFD1 U4693 ( .I(n3930), .Z(n3800) );
  CKBD3 U4694 ( .I(n3931), .Z(n3801) );
  CKBD3 U4695 ( .I(n3869), .Z(n3802) );
  BUFFD2 U4696 ( .I(n3921), .Z(n3803) );
  CKBD3 U4697 ( .I(n3922), .Z(n3804) );
  CKBD3 U4698 ( .I(n3924), .Z(n3805) );
  CKBD3 U4699 ( .I(n3925), .Z(n3806) );
  BUFFD2 U4700 ( .I(n3859), .Z(n3807) );
  CKBD3 U4701 ( .I(n3876), .Z(n3808) );
  CKBD4 U4702 ( .I(n3910), .Z(n3809) );
  CKBD4 U4703 ( .I(n3912), .Z(n3810) );
  CKBD3 U4704 ( .I(n3323), .Z(n3811) );
  CKBD4 U4705 ( .I(n3311), .Z(n3812) );
  BUFFD2 U4706 ( .I(n3721), .Z(n3813) );
  CKBD4 U4707 ( .I(n3673), .Z(n3814) );
  CKBD3 U4708 ( .I(n3674), .Z(n3815) );
  CKBD3 U4709 ( .I(n3675), .Z(n3816) );
  CKBD3 U4710 ( .I(n3676), .Z(n3817) );
  CKBD4 U4711 ( .I(n3724), .Z(n3818) );
  BUFFD2 U4712 ( .I(n3552), .Z(n3819) );
  CKBD3 U4713 ( .I(n3682), .Z(n3820) );
  CKBD3 U4714 ( .I(n3680), .Z(n3821) );
  CKBD3 U4715 ( .I(n3681), .Z(n3822) );
  CKBD3 U4716 ( .I(n3684), .Z(n3823) );
  CKBD3 U4717 ( .I(n3731), .Z(n3824) );
  CKBD3 U4718 ( .I(n3330), .Z(n3825) );
  CKBD3 U4719 ( .I(n3336), .Z(n3826) );
  BUFFD2 U4720 ( .I(n3328), .Z(n3827) );
  BUFFD2 U4721 ( .I(n3335), .Z(n3828) );
  CKBD4 U4722 ( .I(n3703), .Z(n3829) );
  CKBD3 U4723 ( .I(n3505), .Z(n3830) );
  CKBD4 U4724 ( .I(n3750), .Z(n3831) );
  CKBD3 U4725 ( .I(n3865), .Z(n3832) );
  CKBD4 U4726 ( .I(n3872), .Z(n3833) );
  CKBD3 U4727 ( .I(n3671), .Z(n3834) );
  CKBD4 U4728 ( .I(n3672), .Z(n3835) );
  CKBD3 U4729 ( .I(n3669), .Z(n3836) );
  CKBD3 U4730 ( .I(n3666), .Z(n3837) );
  CKBD3 U4731 ( .I(n3667), .Z(n3838) );
  BUFFD1 U4732 ( .I(n3839), .Z(n3128) );
  CKBD1 U4733 ( .I(n3789), .Z(n3977) );
  BUFFD1 U4734 ( .I(n3130), .Z(n3840) );
  BUFFD1 U4735 ( .I(n3909), .Z(n3841) );
  CKBD3 U4736 ( .I(n3916), .Z(n3842) );
  CKBD3 U4737 ( .I(n3920), .Z(n3843) );
  CKBD3 U4738 ( .I(n3923), .Z(n3844) );
  CKBD3 U4739 ( .I(n3960), .Z(n3845) );
  CKBD3 U4740 ( .I(n3962), .Z(n3846) );
  CKBD3 U4741 ( .I(n3963), .Z(n3847) );
  BUFFD1 U4742 ( .I(n3970), .Z(n3848) );
  CKBD3 U4743 ( .I(n3988), .Z(n3849) );
  CKBD3 U4744 ( .I(n3294), .Z(n3850) );
  BUFFD2 U4745 ( .I(n3215), .Z(n3851) );
  CKBD3 U4746 ( .I(n3314), .Z(n3852) );
  CKBD3 U4747 ( .I(n3914), .Z(n3853) );
  CKBD3 U4748 ( .I(n3917), .Z(n3854) );
  CKBD3 U4749 ( .I(n3967), .Z(n3855) );
  CKBD3 U4750 ( .I(n3908), .Z(n3856) );
  CKBD4 U4751 ( .I(n3961), .Z(n3857) );
  CKBD4 U4752 ( .I(n3972), .Z(n3858) );
  BUFFD2 U4753 ( .I(n3313), .Z(n3859) );
  CKBD4 U4754 ( .I(n3331), .Z(n3860) );
  CKBD3 U4755 ( .I(n3719), .Z(n3861) );
  BUFFD2 U4756 ( .I(n3332), .Z(n3862) );
  CKBD4 U4757 ( .I(n3723), .Z(n3863) );
  BUFFD2 U4758 ( .I(n3308), .Z(n3864) );
  CKBD3 U4759 ( .I(n3340), .Z(n3865) );
  CKBD3 U4760 ( .I(n3726), .Z(n3866) );
  BUFFD2 U4761 ( .I(n3334), .Z(n3867) );
  CKBD3 U4762 ( .I(n3338), .Z(n3868) );
  CKBD3 U4763 ( .I(n3339), .Z(n3869) );
  BUFFD2 U4764 ( .I(n3322), .Z(n3870) );
  BUFFD2 U4765 ( .I(n3341), .Z(n3871) );
  CKBD3 U4766 ( .I(n3333), .Z(n3872) );
  CKBD3 U4767 ( .I(n3664), .Z(n3873) );
  BUFFD2 U4768 ( .I(n3140), .Z(n3874) );
  CKBD3 U4769 ( .I(n3918), .Z(n3875) );
  CKBD4 U4770 ( .I(n3773), .Z(n3876) );
  CKBD3 U4771 ( .I(n3716), .Z(n3877) );
  CKBD3 U4772 ( .I(n3717), .Z(n3878) );
  CKBD3 U4773 ( .I(n3670), .Z(n3879) );
  BUFFD2 U4774 ( .I(n3714), .Z(n3880) );
  CKBD4 U4775 ( .I(n3720), .Z(n3881) );
  BUFFD6 U4776 ( .I(n3733), .Z(n3882) );
  BUFFD0 U4777 ( .I(n3128), .Z(n3883) );
  BUFFD2 U4778 ( .I(head[2]), .Z(n3884) );
  BUFFD1 U4779 ( .I(n3792), .Z(n3942) );
  BUFFD2 U4780 ( .I(n2209), .Z(n3885) );
  CKBD4 U4781 ( .I(n4036), .Z(n4010) );
  BUFFD1 U4782 ( .I(n2189), .Z(n3979) );
  BUFFD1 U4783 ( .I(n2192), .Z(n3978) );
  BUFFD1 U4784 ( .I(n4118), .Z(n3886) );
  CKBD3 U4785 ( .I(n2221), .Z(n3887) );
  BUFFD1 U4786 ( .I(n3964), .Z(n3888) );
  BUFFD1 U4787 ( .I(n3966), .Z(n3889) );
  BUFFD1 U4788 ( .I(n3969), .Z(n3890) );
  BUFFD1 U4789 ( .I(n3973), .Z(n3891) );
  CKBD3 U4790 ( .I(n3992), .Z(n3892) );
  CKBD3 U4791 ( .I(n4003), .Z(n3893) );
  BUFFD1 U4792 ( .I(n4016), .Z(n3894) );
  BUFFD1 U4793 ( .I(n4019), .Z(n3895) );
  CKBD3 U4794 ( .I(n3327), .Z(n3896) );
  CKBD3 U4795 ( .I(n4025), .Z(n3897) );
  CKBD3 U4796 ( .I(n4026), .Z(n3898) );
  BUFFD2 U4797 ( .I(n3223), .Z(n3899) );
  BUFFD2 U4798 ( .I(n3218), .Z(n3900) );
  BUFFD2 U4799 ( .I(n3216), .Z(n3901) );
  BUFFD1 U4800 ( .I(n3221), .Z(n3902) );
  CKBD3 U4801 ( .I(n3989), .Z(n3903) );
  CKBD3 U4802 ( .I(n3999), .Z(n3904) );
  CKBD3 U4803 ( .I(n4001), .Z(n3905) );
  CKBD3 U4804 ( .I(n4002), .Z(n3906) );
  BUFFD2 U4805 ( .I(n3309), .Z(n3907) );
  CKBD4 U4806 ( .I(n3820), .Z(n3908) );
  CKBD4 U4807 ( .I(n3818), .Z(n3909) );
  CKBD4 U4808 ( .I(n3316), .Z(n3910) );
  CKBD3 U4809 ( .I(n3317), .Z(n3911) );
  CKBD3 U4810 ( .I(n3779), .Z(n3912) );
  CKBD3 U4811 ( .I(n3776), .Z(n3913) );
  CKBD4 U4812 ( .I(n3330), .Z(n3914) );
  BUFFD2 U4813 ( .I(n3326), .Z(n3915) );
  CKBD3 U4814 ( .I(n3824), .Z(n3916) );
  CKBD4 U4815 ( .I(n3336), .Z(n3917) );
  CKBD3 U4816 ( .I(n3335), .Z(n3918) );
  BUFFD2 U4817 ( .I(n3325), .Z(n3919) );
  BUFFD2 U4818 ( .I(n3725), .Z(n3920) );
  BUFFD2 U4830 ( .I(n3310), .Z(n3921) );
  BUFFD2 U4833 ( .I(n3574), .Z(n3922) );
  BUFFD1 U4849 ( .I(n3328), .Z(n3923) );
  CKBD3 U4850 ( .I(n3337), .Z(n3924) );
  BUFFD2 U4851 ( .I(n3329), .Z(n3925) );
  CKBD3 U4852 ( .I(n3850), .Z(n3926) );
  CKBD4 U4853 ( .I(n3965), .Z(n3927) );
  CKBD3 U4854 ( .I(n3715), .Z(n3928) );
  BUFFD2 U4855 ( .I(n3770), .Z(n3929) );
  CKBD3 U4856 ( .I(n3772), .Z(n3930) );
  CKBD3 U4857 ( .I(n3668), .Z(n3931) );
  CKBD4 U4858 ( .I(n3718), .Z(n3932) );
  CKBD4 U4859 ( .I(n3547), .Z(n3933) );
  BUFFD1 U4860 ( .I(n2276), .Z(n3934) );
  BUFFD1 U4861 ( .I(n2272), .Z(n3935) );
  CKBD1 U4862 ( .I(n2263), .Z(n3983) );
  CKBD1 U4863 ( .I(n3883), .Z(n4006) );
  BUFFD1 U4864 ( .I(n2284), .Z(n3936) );
  BUFFD1 U4865 ( .I(n2288), .Z(n3937) );
  BUFFD1 U4866 ( .I(n2292), .Z(n3938) );
  BUFFD1 U4867 ( .I(n2300), .Z(n3939) );
  BUFFD1 U4868 ( .I(n2197), .Z(n3940) );
  BUFFD1 U4869 ( .I(n2857), .Z(n3941) );
  BUFFD1 U4870 ( .I(n2195), .Z(n3980) );
  CKBD3 U4871 ( .I(n4118), .Z(nextTail_o[0]) );
  CKBD3 U4872 ( .I(n3997), .Z(n3944) );
  BUFFD2 U4873 ( .I(n3996), .Z(n3945) );
  BUFFD1 U4874 ( .I(n2231), .Z(n3946) );
  BUFFD1 U4875 ( .I(n2214), .Z(n3947) );
  BUFFD1 U4876 ( .I(n2234), .Z(n3948) );
  CKBD3 U4877 ( .I(n3994), .Z(n3949) );
  CKBD3 U4878 ( .I(n3995), .Z(n3950) );
  CKBD3 U4879 ( .I(n4004), .Z(n3951) );
  CKBD3 U4880 ( .I(n4017), .Z(n3952) );
  CKBD3 U4881 ( .I(n3990), .Z(n3953) );
  CKBD3 U4882 ( .I(n3991), .Z(n3954) );
  CKBD3 U4883 ( .I(n4000), .Z(n3955) );
  CKBD3 U4884 ( .I(n4020), .Z(n3956) );
  CKBD3 U4885 ( .I(n4021), .Z(n3957) );
  CKBD3 U4886 ( .I(n4023), .Z(n3958) );
  CKBD3 U4887 ( .I(n4024), .Z(n3959) );
  BUFFD2 U4888 ( .I(n3311), .Z(n3960) );
  CKBD3 U4889 ( .I(n3823), .Z(n3961) );
  BUFFD2 U4890 ( .I(n3821), .Z(n3962) );
  BUFFD2 U4891 ( .I(n3822), .Z(n3963) );
  CKBD3 U4892 ( .I(n3338), .Z(n3964) );
  CKBD4 U4893 ( .I(n3873), .Z(n3965) );
  BUFFD2 U4894 ( .I(n3333), .Z(n3966) );
  CKBD4 U4895 ( .I(n3683), .Z(n3967) );
  CKBD4 U4896 ( .I(n3829), .Z(n3968) );
  CKBD3 U4897 ( .I(n3988), .Z(n3969) );
  CKBD3 U4898 ( .I(n3315), .Z(n3970) );
  CKBD4 U4899 ( .I(n3993), .Z(n3971) );
  CKBD3 U4900 ( .I(n3819), .Z(n3972) );
  CKBD3 U4901 ( .I(n3863), .Z(n3973) );
  BUFFD1 U4902 ( .I(n2269), .Z(n3974) );
  BUFFD1 U4903 ( .I(n2859), .Z(n3975) );
  BUFFD1 U4904 ( .I(n2186), .Z(n3976) );
  BUFFD1 U4905 ( .I(completionWriteEn_i), .Z(n3981) );
  BUFFD1 U4906 ( .I(n2244), .Z(n3982) );
  BUFFD1 U4907 ( .I(n3941), .Z(n3984) );
  BUFFD1 U4908 ( .I(n4022), .Z(n3985) );
  BUFFD2 U4909 ( .I(n3217), .Z(n3986) );
  BUFFD1 U4910 ( .I(n2235), .Z(n3987) );
  BUFFD2 U4911 ( .I(n3330), .Z(n3988) );
  CKBD3 U4912 ( .I(n3331), .Z(n3989) );
  CKBD3 U4913 ( .I(n3336), .Z(n3990) );
  CKBD3 U4914 ( .I(n3335), .Z(n3991) );
  BUFFD2 U4915 ( .I(n3866), .Z(n3992) );
  CKBD4 U4916 ( .I(n3926), .Z(n3993) );
  CKBD3 U4917 ( .I(n4025), .Z(n3994) );
  CKBD3 U4918 ( .I(n4026), .Z(n3995) );
  BUFFD2 U4919 ( .I(n3327), .Z(n3996) );
  BUFFD2 U4920 ( .I(n4016), .Z(n3997) );
  CKBD3 U4921 ( .I(n4018), .Z(n3998) );
  BUFFD2 U4922 ( .I(n3322), .Z(n3999) );
  BUFFD2 U4923 ( .I(n3341), .Z(n4000) );
  CKBD3 U4924 ( .I(n3340), .Z(n4001) );
  CKBD3 U4925 ( .I(n3334), .Z(n4002) );
  BUFFD1 U4926 ( .I(n3308), .Z(n4003) );
  CKBD4 U4927 ( .I(n3908), .Z(n4004) );
  BUFFD1 U4928 ( .I(n2179), .Z(n4005) );
  BUFFD0 U4929 ( .I(n2257), .Z(n4007) );
  BUFFD1 U4930 ( .I(n2586), .Z(n4008) );
  BUFFD1 U4931 ( .I(n3884), .Z(n4009) );
  CKBD3 U4932 ( .I(n3242), .Z(n4011) );
  BUFFD2 U4933 ( .I(n3224), .Z(n4012) );
  BUFFD1 U4934 ( .I(n2215), .Z(n4013) );
  BUFFD1 U4935 ( .I(n2245), .Z(n4014) );
  CKBD3 U4936 ( .I(n4037), .Z(n4015) );
  BUFFD2 U4937 ( .I(n3338), .Z(n4016) );
  CKBD3 U4938 ( .I(n3316), .Z(n4017) );
  CKBD3 U4939 ( .I(n3315), .Z(n4018) );
  CKBD3 U4940 ( .I(n3314), .Z(n4019) );
  BUFFD2 U4941 ( .I(n3310), .Z(n4020) );
  CKBD3 U4942 ( .I(n3337), .Z(n4021) );
  BUFFD2 U4943 ( .I(n3326), .Z(n4022) );
  CKBD3 U4944 ( .I(n3319), .Z(n4023) );
  CKBD3 U4945 ( .I(n3325), .Z(n4024) );
  BUFFD2 U4946 ( .I(n3339), .Z(n4025) );
  BUFFD2 U4947 ( .I(n3333), .Z(n4026) );
  BUFFD1 U4948 ( .I(\add_x_6/n1 ), .Z(n4027) );
  BUFFD1 U4949 ( .I(n2182), .Z(n4115) );
  BUFFD1 U4950 ( .I(n2246), .Z(n4028) );
  BUFFD0 U4951 ( .I(n3976), .Z(n4029) );
  BUFFD2 U4952 ( .I(n3884), .Z(n4030) );
  BUFFD1 U4953 ( .I(n4117), .Z(n4031) );
  BUFFD1 U4954 ( .I(n2226), .Z(n4032) );
  BUFFD1 U4955 ( .I(n2219), .Z(n4033) );
  BUFFD1 U4956 ( .I(n2238), .Z(n4034) );
  BUFFD1 U4957 ( .I(n2244), .Z(n4035) );
  BUFFD2 U4958 ( .I(n3703), .Z(n4036) );
  BUFFD2 U4959 ( .I(n3329), .Z(n4037) );
  BUFFD1 U4960 ( .I(n2587), .Z(n4038) );
  CKBD1 U4961 ( .I(n2211), .Z(n4039) );
  BUFFD1 U4962 ( .I(n2239), .Z(n4040) );
  CKBD3 U4963 ( .I(n3240), .Z(n4041) );
  BUFFD2 U4964 ( .I(n2225), .Z(n4116) );
  BUFFD2 U4965 ( .I(n3220), .Z(n4042) );
  BUFFD2 U4966 ( .I(n3222), .Z(n4043) );
  BUFFD2 U4967 ( .I(n3160), .Z(n4044) );
  BUFFD2 U4968 ( .I(n3174), .Z(n4045) );
  BUFFD2 U4969 ( .I(n3173), .Z(n4046) );
  BUFFD2 U4970 ( .I(n3172), .Z(n4047) );
  BUFFD2 U4971 ( .I(n3158), .Z(n4048) );
  BUFFD2 U4972 ( .I(n3157), .Z(n4049) );
  BUFFD1 U4973 ( .I(n3200), .Z(n4050) );
  BUFFD2 U4974 ( .I(n3171), .Z(n4051) );
  BUFFD1 U4975 ( .I(n3199), .Z(n4052) );
  BUFFD2 U4976 ( .I(n3156), .Z(n4053) );
  BUFFD2 U4977 ( .I(n3155), .Z(n4054) );
  BUFFD2 U4978 ( .I(n3154), .Z(n4055) );
  BUFFD2 U4979 ( .I(n3153), .Z(n4056) );
  BUFFD1 U4980 ( .I(n3192), .Z(n4057) );
  BUFFD1 U4981 ( .I(n3191), .Z(n4058) );
  BUFFD1 U4982 ( .I(n3209), .Z(n4059) );
  BUFFD1 U4983 ( .I(n3207), .Z(n4060) );
  BUFFD1 U4984 ( .I(n3189), .Z(n4061) );
  BUFFD1 U4985 ( .I(n3205), .Z(n4062) );
  BUFFD1 U4986 ( .I(n3179), .Z(n4063) );
  BUFFD1 U4987 ( .I(n3206), .Z(n4064) );
  BUFFD1 U4988 ( .I(n3203), .Z(n4065) );
  BUFFD1 U4989 ( .I(n3146), .Z(n4066) );
  BUFFD1 U4990 ( .I(n3193), .Z(n4067) );
  BUFFD1 U4991 ( .I(n3210), .Z(n4068) );
  BUFFD1 U4992 ( .I(n3208), .Z(n4069) );
  BUFFD1 U4993 ( .I(n3194), .Z(n4070) );
  BUFFD1 U4994 ( .I(n3204), .Z(n4071) );
  BUFFD1 U4995 ( .I(n3177), .Z(n4072) );
  BUFFD1 U4996 ( .I(n3202), .Z(n4073) );
  BUFFD1 U4997 ( .I(n3196), .Z(n4074) );
  BUFFD1 U4998 ( .I(n3141), .Z(n4075) );
  BUFFD1 U4999 ( .I(n3187), .Z(n4076) );
  BUFFD2 U5000 ( .I(n3178), .Z(n4077) );
  BUFFD1 U5001 ( .I(n3201), .Z(n4078) );
  BUFFD1 U5002 ( .I(n3143), .Z(n4079) );
  BUFFD1 U5003 ( .I(n3145), .Z(n4080) );
  BUFFD2 U5004 ( .I(n3180), .Z(n4081) );
  BUFFD1 U5005 ( .I(n3197), .Z(n4082) );
  BUFFD1 U5006 ( .I(n3142), .Z(n4083) );
  BUFFD1 U5007 ( .I(n3149), .Z(n4084) );
  BUFFD1 U5008 ( .I(n3195), .Z(n4085) );
  BUFFD1 U5009 ( .I(n3198), .Z(n4086) );
  BUFFD1 U5010 ( .I(n3150), .Z(n4087) );
  BUFFD1 U5011 ( .I(n3144), .Z(n4088) );
  BUFFD1 U5012 ( .I(n3147), .Z(n4089) );
  BUFFD2 U5013 ( .I(n3148), .Z(n4090) );
  BUFFD2 U5014 ( .I(n3151), .Z(n4091) );
  BUFFD1 U5015 ( .I(n3163), .Z(n4092) );
  BUFFD1 U5016 ( .I(n3164), .Z(n4093) );
  BUFFD2 U5017 ( .I(n3186), .Z(n4094) );
  BUFFD2 U5018 ( .I(n3183), .Z(n4095) );
  BUFFD2 U5019 ( .I(n3219), .Z(n4096) );
  BUFFD2 U5020 ( .I(n3182), .Z(n4097) );
  BUFFD2 U5021 ( .I(n3165), .Z(n4098) );
  BUFFD1 U5022 ( .I(n3152), .Z(n4099) );
  BUFFD2 U5023 ( .I(n3184), .Z(n4100) );
  BUFFD2 U5024 ( .I(n3181), .Z(n4101) );
  BUFFD2 U5025 ( .I(n3190), .Z(n4102) );
  BUFFD2 U5026 ( .I(n3169), .Z(n4103) );
  BUFFD2 U5027 ( .I(n3175), .Z(n4104) );
  BUFFD2 U5028 ( .I(n3170), .Z(n4105) );
  BUFFD2 U5029 ( .I(n3176), .Z(n4106) );
  BUFFD2 U5030 ( .I(n3188), .Z(n4107) );
  BUFFD2 U5031 ( .I(n3185), .Z(n4108) );
  BUFFD2 U5032 ( .I(n3168), .Z(n4109) );
  BUFFD2 U5033 ( .I(n3167), .Z(n4110) );
  BUFFD2 U5034 ( .I(n3166), .Z(n4111) );
  BUFFD2 U5035 ( .I(n3162), .Z(n4112) );
  BUFFD2 U5036 ( .I(n3161), .Z(n4113) );
  BUFFD2 U5037 ( .I(n3159), .Z(n4114) );
  BUFFD2 U5038 ( .I(reset_i), .Z(n4117) );
endmodule

