library verilog;
use verilog.vl_types.all;
entity divider_testbench is
end divider_testbench;
