../../src/verilog/forwardingUnit.sv