../../src/verilog/instructionFetch.sv