../../src/verilog/orGate16.sv