../../src/verilog/signExtend9.sv