../../src/verilog/registerX16.sv