library verilog;
use verilog.vl_types.all;
entity mux4x1_testbench is
end mux4x1_testbench;
