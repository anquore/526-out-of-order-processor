../../src/verilog/norifier.sv