library verilog;
use verilog.vl_types.all;
entity orGate16_testbench is
end orGate16_testbench;
