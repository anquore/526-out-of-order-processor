../../src/verilog/decoder1x2.sv