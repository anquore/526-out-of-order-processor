../../src/syn/netlist/ROB.sv