../../src/verilog/NAND_MUX_4x1.sv