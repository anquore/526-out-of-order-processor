../../src/verilog/datamem.sv