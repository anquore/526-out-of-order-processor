library verilog;
use verilog.vl_types.all;
entity decodeStage_testbench is
end decodeStage_testbench;
