library verilog;
use verilog.vl_types.all;
entity bitSlice_testbench is
end bitSlice_testbench;
