../../src/verilog/ROBregs.sv