../../src/verilog/shiftLeft2.sv