../../src/verilog/registerX64.sv