library verilog;
use verilog.vl_types.all;
entity NAND_MUX_4x1_testbench is
end NAND_MUX_4x1_testbench;
