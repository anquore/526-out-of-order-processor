library verilog;
use verilog.vl_types.all;
entity NAND_MUX_2x1_testbench is
end NAND_MUX_2x1_testbench;
