../../src/verilog/fullAdder.sv