../../src/verilog/memStage.sv