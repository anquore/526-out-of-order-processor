../../src/verilog/pipelined.sv