../../src/verilog/mux_2x1_X64.sv