../../src/verilog/instructmem.sv