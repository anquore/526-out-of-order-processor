../../src/verilog/mux16x1.sv