../../src/verilog/signExtend26.sv