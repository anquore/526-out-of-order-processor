../../src/verilog/divider.sv