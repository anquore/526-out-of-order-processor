library verilog;
use verilog.vl_types.all;
entity mux2x5_testbench is
end mux2x5_testbench;
