../../src/verilog/control.sv