../../src/verilog/full_adder.sv