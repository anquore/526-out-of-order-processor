../../src/verilog/FF_en.sv