library verilog;
use verilog.vl_types.all;
entity adder64_testbench is
end adder64_testbench;
